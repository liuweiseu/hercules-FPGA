.box 1 mipi_rx_pinf_tx_pinf_1080_ipc_adder_12 25 13
.input 1 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11]
.output 1 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11]
.delay 1
1300	1200	1100	1000	900	800	700	600	500	400	300	200	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 2 mipi_rx_pinf_tx_pinf_1080_ipc_adder_9 19 10
.input 2 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8]
.output 2 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8]
.delay 2
1000	900	800	700	600	500	400	300	200	900	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	500	600	500	400	300	200	-	-	-	-	
700	600	500	400	300	200	-	-	-	600	700	600	500	400	300	200	-	-	-	
800	700	600	500	400	300	200	-	-	700	800	700	600	500	400	300	200	-	-	
900	800	700	600	500	400	300	200	-	800	900	800	700	600	500	400	300	200	-	
1000	900	800	700	600	500	400	300	200	900	1000	900	800	700	600	500	400	300	200	


.box 3 mipi_rx_pinf_tx_pinf_1080_ipc_adder_13 27 14
.input 3 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12]
.output 3 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12]
.delay 3
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 4 mipi_rx_pinf_tx_pinf_1080_ipc_adder_11 23 12
.input 4 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10]
.output 4 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10]
.delay 4
1200	1100	1000	900	800	700	600	500	400	300	200	1100	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	
1200	1100	1000	900	800	700	600	500	400	300	200	1100	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 5 mipi_rx_pinf_tx_pinf_1080_ipc_adder_8 17 9
.input 5 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7]
.output 5 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7]
.delay 5
900	800	700	600	500	400	300	200	800	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	300	400	300	200	-	-	-	-	-	
500	400	300	200	-	-	-	-	400	500	400	300	200	-	-	-	-	
600	500	400	300	200	-	-	-	500	600	500	400	300	200	-	-	-	
700	600	500	400	300	200	-	-	600	700	600	500	400	300	200	-	-	
800	700	600	500	400	300	200	-	700	800	700	600	500	400	300	200	-	
900	800	700	600	500	400	300	200	800	900	800	700	600	500	400	300	200	


