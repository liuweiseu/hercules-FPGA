//2018-09-18 glliu
//Add simulation model of H6_BASIC_IO, H6_IOC_FUN.

`timescale 1ns/1ps
//----------------------------------------------------------------------------
//
// module: ADD1_A
//
// description:     1-bit full adder with invertable a input
//
//----------------------------------------------------------------------------

module ADD1_A (
        a,
        b,
        ci,
        co,
        s
        );
        
    input       a;
    input       b;
    input       ci;
    output      co;
    output      s;
    
    parameter a_inv = "false";   //a input invert, default is "false"

    wire a_in;
    assign a_in = (a_inv == "false") ?  a : ~a;
    assign p  = a_in ^ b;
    assign pb = ~p;
    assign co = p ? ci : a_in ;
    assign s  = ci ^ p;

endmodule



module GND (Y);
    output Y;
    
    assign Y = 0;

endmodule


//----------------------------------------------------------------------------
//
// module: IBUF
//
// description:     input buffer
//
//----------------------------------------------------------------------------

module IBUF (p, o);
    input   p;
    output  o;

    buf b1 (o, p);

endmodule

//----------------------------------------------------------------------------
//
// module: IOBUF
//
// description:     Multiplexer of IOCLK 
//
//----------------------------------------------------------------------------
module IOBUF(
    i0,
    i1,
    i2,
    i3,
    i4,
    i5,
    i6,
    i7,
    o
);

input           i0;
input           i1;
input           i2;
input           i3;
input           i4;
input           i5;
input           i6;
input           i7;
output          o;

parameter SEL = 6'b00000;

wire Z0,Z1;
assign   Z0 =
              (SEL[3:0] == 4'b0001) ? i0 :
              (SEL[3:0] == 4'b0010) ? i1 :
              (SEL[3:0] == 4'b0100) ? i2 : 
              (SEL[3:0] == 4'b1000) ? i3 : 
              (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
assign   Z1 =
              (SEL[3:0] == 4'b0001) ? i4 :
              (SEL[3:0] == 4'b0010) ? i5 :
              (SEL[3:0] == 4'b0100) ? i6 : 
              (SEL[3:0] == 4'b1000) ? i7 : 
              (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
assign	 o =
              (SEL[5:4] == 2'b01) ? Z0 :
              (SEL[5:4] == 2'b10) ? Z1 :
              (SEL[5:4] == 2'b00) ? 1'b0 : 1'bx;

endmodule

module IOC (
    id,
    od,
    clk,
    rstn,
    setn,
    clk_en,
    oen,
    pad 
);

    output        id;     //output data to fabric
    input        od;     //input data from fabric
    input        oen;
    input       clk;
    input       clk_en;
    input       rstn;
    input       setn;
    inout        pad;
    

    parameter slew_rate = "fastest";//slowest,slow,fast,fastest
    parameter driving_strength = "16ma";//base,4ma,8ma,12ma,16ma
    parameter keep_sel = "none";//pullup,keep,none,pulldown
    
    parameter reg_always_en = "false";  //true, false
    parameter is_en_used = "false";     //true, false

    parameter is_rstn_inv = "false";    //true
    parameter is_setn_inv = "false";    //true
    parameter is_clk_inv  = "false";    //true
    parameter is_od_inv = "false";      //true
    parameter is_oen_inv = "false";     //true

    parameter oen_sel = "vcc";        //register, gnd(output), vcc(input)
    parameter od_sel = "gnd";         //register, gnd, vcc,bypass
    parameter id_sel = "bypass";      //register
    
    parameter oen_setn_en = "false"; //true
    parameter oen_rstn_en = "false"; //true

    parameter od_setn_en = "false"; //true
    parameter od_rstn_en = "false"; //true
    
    parameter id_setn_en = "false"; //true
    parameter id_rstn_en = "false"; //true

    parameter optional_function = ""; //"spi_sclk", "spi_sdi", "spi_cson", "spi_sdo", ""
    
    wire i_clk;
    wire i_rstn;
    wire i_setn;
    wire i_oen;
    wire i_od;
    
    wire     id_reg;
    wire    od_reg;
    wire    oen_reg;

    wire    id_rstn;
    wire    id_setn;
    wire    od_rstn;
    wire    od_setn;
    wire    oen_setn;
    wire    oen_rstn;

    wire    en;
    wire    out_en;
    wire    out_data;

    
    /*---------- inverted setting----------------*/      
    assign i_clk    = (is_clk_inv  == "true") ? ~clk : clk;      
    assign i_oen    = (is_oen_inv  == "true") ? ~oen : oen;       
    assign i_od     = (is_od_inv   == "true") ? ~od : od;       
    assign en       = (reg_always_en == "true") ? 1'b1 : (is_en_used == "true" ? clk_en : 1'b0);
    assign i_rstn   = (is_rstn_inv == "true") ? ~rstn : rstn;       
    assign i_setn   = (is_setn_inv == "true") ? ~setn : setn;       

    assign id_rstn  = (id_rstn_en == "true") ? i_rstn : 1'b1;
    assign id_setn  = (id_setn_en == "true") ? i_setn : 1'b1;

    assign od_rstn  = (od_rstn_en == "true") ? i_rstn : 1'b1;
    assign od_setn  = (od_setn_en == "true") ? i_setn : 1'b1;

    assign oen_rstn  = (oen_rstn_en == "true") ? i_rstn : 1'b1;
    assign oen_setn  = (oen_setn_en == "true") ? i_setn : 1'b1;

    /*---------- id Reg----------------*/  
    DFFRSEN IPREGDFF(.Q (id_reg), .D (pad), .CLK (i_clk), .RST (~id_rstn), .SET(~id_setn), .EN(en));
    
    /*---------- od Reg----------------*/  
    DFFRSEN OPREGDFF(.Q (od_reg), .D (i_od), .CLK (i_clk), .RST (~od_rstn), .SET(~od_setn), .EN(en));

    /*---------- Oe Reg----------------*/  
    DFFRSEN OEPREGDFF(.Q (oen_reg), .D (i_oen), .CLK (i_clk), .RST (~oen_rstn), .SET(~oen_setn), .EN(en));
    
    /*---------- Input Generation----------------*/
    assign id = (id_sel == "register") ? id_reg : pad;
    
    /*---------- Oen Generation----------------*/
    assign out_en = (oen_sel == "register") ? oen_reg :
                    (oen_sel == "bypass")   ? i_oen :
                    (oen_sel == "vcc")  ? 1'b1 :
                    (oen_sel == "gnd")  ? 1'b0 : 1'bx;
                                    
    /*---------- Output Generation----------------*/
    assign out_data = (od_sel == "register") ? od_reg :
                      (od_sel == "bypass" )  ? i_od :
                      (od_sel == "vcc") ? 1'b1 :
                      (od_sel == "gnd") ? 1'b0 : 1'bx;

    assign pad = ~out_en ? out_data : 1'bz;


endmodule

module DFFRSEN (Q, D, CLK, RST, SET, EN);
    input    D;
    input    CLK;
    input    EN;
    input    RST;
    input    SET;
    output    Q;
    
    reg        qo;
    
    always @(posedge CLK or posedge RST or posedge SET)
        if(RST)
            qo <= 1'b0;
        else if (SET)
            qo <= 1'b1;
        else if(EN)
            qo <= D;
    
    assign Q = qo;
    
endmodule


//----------------------------------------------------------------------------
//
// module: LUT5_2
//
// description: 5 input, 2 outputs lookup-table
// config_x:      32 bit init value
// config_y:      32 bit init value
//
//----------------------------------------------------------------------------

module LUT5_2 (
         dx,
         dy,
         f4,
         f3,
         f2,
         f1,
         f0
         );

    input       f4;
    input       f3;
    input       f2;
    input       f1;
    input       f0;

    output      dx;
    output      dy;

    parameter       config_data_x = 32'h0000_0000;
    parameter       config_data_y = 32'h0000_0000;

    wire [31:0]         cfg_x = config_data_x;
    wire [31:0]         cfg_xy = config_data_y;
      
    wire [15:0]         da_x;
    wire [7:0]          db_x;
    wire [3:0]          dc_x;
    wire [1:0]          dd_x;
    wire                de_x;

    wire [15:0]         da_xy;
    wire [7:0]          db_xy;
    wire [3:0]          dc_xy;
    wire [1:0]          dd_xy;
    wire                de_xy;
    //LUT5_X
    MUX2S_L muxa0_x(.o(da_x[0]),  .sel(f0), .i1(cfg_x[1]), .i0(cfg_x[0]) );
    MUX2S_L muxa1_x(.o(da_x[1]),  .sel(f0), .i1(cfg_x[3]), .i0(cfg_x[2]) );
    MUX2S_L muxa2_x(.o(da_x[2]),  .sel(f0), .i1(cfg_x[5]), .i0(cfg_x[4]) );
    MUX2S_L muxa3_x(.o(da_x[3]),  .sel(f0), .i1(cfg_x[7]), .i0(cfg_x[6]) );
    MUX2S_L muxa4_x(.o(da_x[4]),  .sel(f0), .i1(cfg_x[9]), .i0(cfg_x[8]) );
    MUX2S_L muxa5_x(.o(da_x[5]),  .sel(f0), .i1(cfg_x[11]), .i0(cfg_x[10]) );
    MUX2S_L muxa6_x(.o(da_x[6]),  .sel(f0), .i1(cfg_x[13]), .i0(cfg_x[12]) );
    MUX2S_L muxa7_x(.o(da_x[7]),  .sel(f0), .i1(cfg_x[15]), .i0(cfg_x[14]) );
    MUX2S_L muxa8_x(.o(da_x[8]),  .sel(f0), .i1(cfg_x[17]), .i0(cfg_x[16]) );
    MUX2S_L muxa9_x(.o(da_x[9]),  .sel(f0), .i1(cfg_x[19]), .i0(cfg_x[18]) );
    MUX2S_L muxa10_x(.o(da_x[10]), .sel(f0), .i1(cfg_x[21]), .i0(cfg_x[20]) );
    MUX2S_L muxa11_x(.o(da_x[11]), .sel(f0), .i1(cfg_x[23]), .i0(cfg_x[22]) );
    MUX2S_L muxa12_x(.o(da_x[12]), .sel(f0), .i1(cfg_x[25]), .i0(cfg_x[24]) );
    MUX2S_L muxa13_x(.o(da_x[13]), .sel(f0), .i1(cfg_x[27]), .i0(cfg_x[26]) );
    MUX2S_L muxa14_x(.o(da_x[14]), .sel(f0), .i1(cfg_x[29]), .i0(cfg_x[28]) );
    MUX2S_L muxa15_x(.o(da_x[15]), .sel(f0), .i1(cfg_x[31]), .i0(cfg_x[30]) );

    MUX2S_L muxb0_x(.o(db_x[0]), .sel(f1), .i1(da_x[1]), .i0(da_x[0]) );
    MUX2S_L muxb1_x(.o(db_x[1]), .sel(f1), .i1(da_x[3]), .i0(da_x[2]) );
    MUX2S_L muxb2_x(.o(db_x[2]), .sel(f1), .i1(da_x[5]), .i0(da_x[4]) );
    MUX2S_L muxb3_x(.o(db_x[3]), .sel(f1), .i1(da_x[7]), .i0(da_x[6]) );
    MUX2S_L muxb4_x(.o(db_x[4]), .sel(f1), .i1(da_x[9]), .i0(da_x[8]) );
    MUX2S_L muxb5_x(.o(db_x[5]), .sel(f1), .i1(da_x[11]), .i0(da_x[10]) );
    MUX2S_L muxb6_x(.o(db_x[6]), .sel(f1), .i1(da_x[13]), .i0(da_x[12]) );
    MUX2S_L muxb7_x(.o(db_x[7]), .sel(f1), .i1(da_x[15]), .i0(da_x[14]) );

    MUX2S_L muxc0_x(.o(dc_x[0]), .sel(f2), .i1(db_x[1]), .i0(db_x[0]) );
    MUX2S_L muxc1_x(.o(dc_x[1]), .sel(f2), .i1(db_x[3]), .i0(db_x[2]) );
    MUX2S_L muxc2_x(.o(dc_x[2]), .sel(f2), .i1(db_x[5]), .i0(db_x[4]) );
    MUX2S_L muxc3_x(.o(dc_x[3]), .sel(f2), .i1(db_x[7]), .i0(db_x[6]) );

    MUX2S_L muxd0_x(.o(dd_x[0]), .sel(f3), .i1(dc_x[1]), .i0(dc_x[0]) );
    MUX2S_L muxd1_x(.o(dd_x[1]), .sel(f3), .i1(dc_x[3]), .i0(dc_x[2]) );

    MUX2S_L muxe0_x(.o(de_x), .sel(f4), .i1(dd_x[1]), .i0(dd_x[0]) );

    //LUT5_XY
    MUX2S_L muxa0_xy(.o(da_xy[0]),  .sel(f0), .i1(cfg_xy[1]), .i0(cfg_xy[0]) );
    MUX2S_L muxa1_xy(.o(da_xy[1]),  .sel(f0), .i1(cfg_xy[3]), .i0(cfg_xy[2]) );
    MUX2S_L muxa2_xy(.o(da_xy[2]),  .sel(f0), .i1(cfg_xy[5]), .i0(cfg_xy[4]) );
    MUX2S_L muxa3_xy(.o(da_xy[3]),  .sel(f0), .i1(cfg_xy[7]), .i0(cfg_xy[6]) );
    MUX2S_L muxa4_xy(.o(da_xy[4]),  .sel(f0), .i1(cfg_xy[9]), .i0(cfg_xy[8]) );
    MUX2S_L muxa5_xy(.o(da_xy[5]),  .sel(f0), .i1(cfg_xy[11]), .i0(cfg_xy[10]) );
    MUX2S_L muxa6_xy(.o(da_xy[6]),  .sel(f0), .i1(cfg_xy[13]), .i0(cfg_xy[12]) );
    MUX2S_L muxa7_xy(.o(da_xy[7]),  .sel(f0), .i1(cfg_xy[15]), .i0(cfg_xy[14]) );
    MUX2S_L muxa8_xy(.o(da_xy[8]),  .sel(f0), .i1(cfg_xy[17]), .i0(cfg_xy[16]) );
    MUX2S_L muxa9_xy(.o(da_xy[9]),  .sel(f0), .i1(cfg_xy[19]), .i0(cfg_xy[18]) );
    MUX2S_L muxa10_xy(.o(da_xy[10]), .sel(f0), .i1(cfg_xy[21]), .i0(cfg_xy[20]) );
    MUX2S_L muxa11_xy(.o(da_xy[11]), .sel(f0), .i1(cfg_xy[23]), .i0(cfg_xy[22]) );
    MUX2S_L muxa12_xy(.o(da_xy[12]), .sel(f0), .i1(cfg_xy[25]), .i0(cfg_xy[24]) );
    MUX2S_L muxa13_xy(.o(da_xy[13]), .sel(f0), .i1(cfg_xy[27]), .i0(cfg_xy[26]) );
    MUX2S_L muxa14_xy(.o(da_xy[14]), .sel(f0), .i1(cfg_xy[29]), .i0(cfg_xy[28]) );
    MUX2S_L muxa15_xy(.o(da_xy[15]), .sel(f0), .i1(cfg_xy[31]), .i0(cfg_xy[30]) );

    MUX2S_L muxb0_xy(.o(db_xy[0]), .sel(f1), .i1(da_xy[1]), .i0(da_xy[0]) );
    MUX2S_L muxb1_xy(.o(db_xy[1]), .sel(f1), .i1(da_xy[3]), .i0(da_xy[2]) );
    MUX2S_L muxb2_xy(.o(db_xy[2]), .sel(f1), .i1(da_xy[5]), .i0(da_xy[4]) );
    MUX2S_L muxb3_xy(.o(db_xy[3]), .sel(f1), .i1(da_xy[7]), .i0(da_xy[6]) );
    MUX2S_L muxb4_xy(.o(db_xy[4]), .sel(f1), .i1(da_xy[9]), .i0(da_xy[8]) );
    MUX2S_L muxb5_xy(.o(db_xy[5]), .sel(f1), .i1(da_xy[11]), .i0(da_xy[10]) );
    MUX2S_L muxb6_xy(.o(db_xy[6]), .sel(f1), .i1(da_xy[13]), .i0(da_xy[12]) );
    MUX2S_L muxb7_xy(.o(db_xy[7]), .sel(f1), .i1(da_xy[15]), .i0(da_xy[14]) );

    MUX2S_L muxc0_xy(.o(dc_xy[0]), .sel(f2), .i1(db_xy[1]), .i0(db_xy[0]) );
    MUX2S_L muxc1_xy(.o(dc_xy[1]), .sel(f2), .i1(db_xy[3]), .i0(db_xy[2]) );
    MUX2S_L muxc2_xy(.o(dc_xy[2]), .sel(f2), .i1(db_xy[5]), .i0(db_xy[4]) );
    MUX2S_L muxc3_xy(.o(dc_xy[3]), .sel(f2), .i1(db_xy[7]), .i0(db_xy[6]) );

    MUX2S_L muxd0_xy(.o(dd_xy[0]), .sel(f3), .i1(dc_xy[1]), .i0(dc_xy[0]) );
    MUX2S_L muxd1_xy(.o(dd_xy[1]), .sel(f3), .i1(dc_xy[3]), .i0(dc_xy[2]) );

    MUX2S_L muxe0_xy(.o(de_xy), .sel(f4), .i1(dd_xy[1]), .i0(dd_xy[0]) );

    assign        dx = de_x;
    assign        dy = de_xy;

endmodule


//----------------------------------------------------------------------------
//
// module: LUT6
//
// description: 6 input lookup-table
// config:      64 bit init value
//
//----------------------------------------------------------------------------

module LUT6 (
         xy,
         f5,
         f4,
         f3,
         f2,
         f1,
         f0
         );

    input       f5;
    input       f4;
    input       f3;
    input       f2;
    input       f1;
    input       f0;

    output      xy;

    parameter       config_data = 64'h0000_0000_0000_0000;

    wire [63:0]         cfg = config_data;
    wire [31:0]         da;
    wire [15:0]         db;
    wire [7:0]          dc;
    wire [3:0]          dd;
    wire [1:0]          de;
    wire                df;

    MUX2S_L muxa0 (.o(da[0]),  .sel(f0), .i1(cfg[1]),  .i0(cfg[0]) );
    MUX2S_L muxa1 (.o(da[1]),  .sel(f0), .i1(cfg[3]),  .i0(cfg[2]) );
    MUX2S_L muxa2 (.o(da[2]),  .sel(f0), .i1(cfg[5]),  .i0(cfg[4]) );
    MUX2S_L muxa3 (.o(da[3]),  .sel(f0), .i1(cfg[7]),  .i0(cfg[6]) );
    MUX2S_L muxa4 (.o(da[4]),  .sel(f0), .i1(cfg[9]),  .i0(cfg[8]) );
    MUX2S_L muxa5 (.o(da[5]),  .sel(f0), .i1(cfg[11]), .i0(cfg[10]) );
    MUX2S_L muxa6 (.o(da[6]),  .sel(f0), .i1(cfg[13]), .i0(cfg[12]) );
    MUX2S_L muxa7 (.o(da[7]),  .sel(f0), .i1(cfg[15]), .i0(cfg[14]) );
    MUX2S_L muxa8 (.o(da[8]),  .sel(f0), .i1(cfg[17]), .i0(cfg[16]) );
    MUX2S_L muxa9 (.o(da[9]),  .sel(f0), .i1(cfg[19]), .i0(cfg[18]) );
    MUX2S_L muxa10(.o(da[10]), .sel(f0), .i1(cfg[21]), .i0(cfg[20]) );
    MUX2S_L muxa11(.o(da[11]), .sel(f0), .i1(cfg[23]), .i0(cfg[22]) );
    MUX2S_L muxa12(.o(da[12]), .sel(f0), .i1(cfg[25]), .i0(cfg[24]) );
    MUX2S_L muxa13(.o(da[13]), .sel(f0), .i1(cfg[27]), .i0(cfg[26]) );
    MUX2S_L muxa14(.o(da[14]), .sel(f0), .i1(cfg[29]), .i0(cfg[28]) );
    MUX2S_L muxa15(.o(da[15]), .sel(f0), .i1(cfg[31]), .i0(cfg[30]) );
    MUX2S_L muxa16(.o(da[16]), .sel(f0), .i1(cfg[33]), .i0(cfg[32]) );
    MUX2S_L muxa17(.o(da[17]), .sel(f0), .i1(cfg[35]), .i0(cfg[34]) );
    MUX2S_L muxa18(.o(da[18]), .sel(f0), .i1(cfg[37]), .i0(cfg[36]) );
    MUX2S_L muxa19(.o(da[19]), .sel(f0), .i1(cfg[39]), .i0(cfg[38]) );
    MUX2S_L muxa20(.o(da[20]), .sel(f0), .i1(cfg[41]), .i0(cfg[40]) );
    MUX2S_L muxa21(.o(da[21]), .sel(f0), .i1(cfg[43]), .i0(cfg[42]) );
    MUX2S_L muxa22(.o(da[22]), .sel(f0), .i1(cfg[45]), .i0(cfg[44]) );
    MUX2S_L muxa23(.o(da[23]), .sel(f0), .i1(cfg[47]), .i0(cfg[46]) );
    MUX2S_L muxa24(.o(da[24]), .sel(f0), .i1(cfg[49]), .i0(cfg[48]) );
    MUX2S_L muxa25(.o(da[25]), .sel(f0), .i1(cfg[51]), .i0(cfg[50]) );
    MUX2S_L muxa26(.o(da[26]), .sel(f0), .i1(cfg[53]), .i0(cfg[52]) );
    MUX2S_L muxa27(.o(da[27]), .sel(f0), .i1(cfg[55]), .i0(cfg[54]) );
    MUX2S_L muxa28(.o(da[28]), .sel(f0), .i1(cfg[57]), .i0(cfg[56]) );
    MUX2S_L muxa29(.o(da[29]), .sel(f0), .i1(cfg[59]), .i0(cfg[58]) );
    MUX2S_L muxa30(.o(da[30]), .sel(f0), .i1(cfg[61]), .i0(cfg[60]) );
    MUX2S_L muxa31(.o(da[31]), .sel(f0), .i1(cfg[63]), .i0(cfg[62]) );

    MUX2S_L muxb0 (.o(db[0]),  .sel(f1), .i1(da[1]),  .i0(da[0]) );
    MUX2S_L muxb1 (.o(db[1]),  .sel(f1), .i1(da[3]),  .i0(da[2]) );
    MUX2S_L muxb2 (.o(db[2]),  .sel(f1), .i1(da[5]),  .i0(da[4]) );
    MUX2S_L muxb3 (.o(db[3]),  .sel(f1), .i1(da[7]),  .i0(da[6]) );
    MUX2S_L muxb4 (.o(db[4]),  .sel(f1), .i1(da[9]),  .i0(da[8]) );
    MUX2S_L muxb5 (.o(db[5]),  .sel(f1), .i1(da[11]), .i0(da[10]) );
    MUX2S_L muxb6 (.o(db[6]),  .sel(f1), .i1(da[13]), .i0(da[12]) );
    MUX2S_L muxb7 (.o(db[7]),  .sel(f1), .i1(da[15]), .i0(da[14]) );
    MUX2S_L muxb8 (.o(db[8]),  .sel(f1), .i1(da[17]), .i0(da[16]) );
    MUX2S_L muxb9 (.o(db[9]),  .sel(f1), .i1(da[19]), .i0(da[18]) );
    MUX2S_L muxb10(.o(db[10]), .sel(f1), .i1(da[21]), .i0(da[20]) );
    MUX2S_L muxb11(.o(db[11]), .sel(f1), .i1(da[23]), .i0(da[22]) );
    MUX2S_L muxb12(.o(db[12]), .sel(f1), .i1(da[25]), .i0(da[24]) );
    MUX2S_L muxb13(.o(db[13]), .sel(f1), .i1(da[27]), .i0(da[26]) );
    MUX2S_L muxb14(.o(db[14]), .sel(f1), .i1(da[29]), .i0(da[28]) );
    MUX2S_L muxb15(.o(db[15]), .sel(f1), .i1(da[31]), .i0(da[30]) );

    MUX2S_L muxc0(.o(dc[0]), .sel(f2), .i1(db[1]),  .i0(db[0]) );
    MUX2S_L muxc1(.o(dc[1]), .sel(f2), .i1(db[3]),  .i0(db[2]) );
    MUX2S_L muxc2(.o(dc[2]), .sel(f2), .i1(db[5]),  .i0(db[4]) );
    MUX2S_L muxc3(.o(dc[3]), .sel(f2), .i1(db[7]),  .i0(db[6]) );
    MUX2S_L muxc4(.o(dc[4]), .sel(f2), .i1(db[9]),  .i0(db[8]) );
    MUX2S_L muxc5(.o(dc[5]), .sel(f2), .i1(db[11]), .i0(db[10]) );
    MUX2S_L muxc6(.o(dc[6]), .sel(f2), .i1(db[13]), .i0(db[12]) );
    MUX2S_L muxc7(.o(dc[7]), .sel(f2), .i1(db[15]), .i0(db[14]) );

    MUX2S_L muxd0(.o(dd[0]), .sel(f3), .i1(dc[1]), .i0(dc[0]) );
    MUX2S_L muxd1(.o(dd[1]), .sel(f3), .i1(dc[3]), .i0(dc[2]) );
    MUX2S_L muxd2(.o(dd[2]), .sel(f3), .i1(dc[5]), .i0(dc[4]) );
    MUX2S_L muxd3(.o(dd[3]), .sel(f3), .i1(dc[7]), .i0(dc[6]) );

    MUX2S_L muxe0(.o(de[0]), .sel(f4), .i1(dd[1]), .i0(dd[0]) );
    MUX2S_L muxe1(.o(de[1]), .sel(f4), .i1(dd[3]), .i0(dd[2]) );

    MUX2S_L muxf0(.o(df), .sel(f5), .i1(de[1]), .i0(de[0]) );

    assign      xy = df;

endmodule

//----------------------------------------------------------------------------
//
// module: MUXF7
//
// description:     2-to-1 MUXF7 
//
//----------------------------------------------------------------------------

module MUXF7 (
          out,
          sel,
          in0,
          in1
          );

   input        in0;
   input        in1;
   input        sel;

   output       out; 

   assign       out = (sel == 1'b0) ? in0 :
                      (sel == 1'b1) ? in1 : 1'bx;

endmodule


//----------------------------------------------------------------------------
//
// module: MUXF8
//
// description:     2-to-1 MUXF8
//
//----------------------------------------------------------------------------

module MUXF8 (
          out,
          sel,
          in0,
          in1
          );

   input        in0;
   input        in1;
   input        sel;

   output       out; 

   assign       out = (sel == 1'b0) ? in0 :
                      (sel == 1'b1) ? in1 : 1'bx;

endmodule


//----------------------------------------------------------------------------
//
// module: OBUF
//
// description:     output buffer
//
//----------------------------------------------------------------------------

module OBUF (p, i);
    input   i;
    output  p;

    buf b1 (p, i);

endmodule


//----------------------------------------------------------------------------
//
// module: OBUFT
//
// description:     tri-state output buffer
//
//----------------------------------------------------------------------------

module OBUFT (p, i, oe);
    input   i;
    input   oe;
    output  p;
    
    bufif0 t1 (p, i, oe);
   
endmodule


//----------------------------------------------------------------------------
//
// module: REG
//
// description:     1-bit register 
//
//----------------------------------------------------------------------------

module REG (
    qx ,
    di ,
    sr ,
    en ,
    clk 
);

parameter   init            = 1'b0;     //register initial value, default is "1'b0"
parameter   sr_value        = 1'b0;     //output value of reset, default is "1'b0"


parameter   always_en       = 1'b0;     //0 for use external enable, 1 for always enable, default is "1'b0"
parameter   no_sr           = 1'b0;     //0 for use external set/reset, 1 for no set/reset, default is "1'b0"
parameter   latch_mode      = 1'b0;     //0 for register mode, 1 for latch mode, default is "1'b0"
parameter   sync_mode       = 1'b0;     //0 for asynchronous mode, 1 for synchronous mode, default is "1'b0"
parameter   clk_inv         = 1'b0;     //0 for clock not inverted, 1 for clock inverted, default is "1'b0"
parameter   en_inv          = 1'b0;     //0 for enable not inverted, 1 for enable inverted, default is "1'b0"
parameter   sr_inv          = 1'b0;     //0 for sr not inverted, 1 for sr inverted, default is "1'b0"

output  qx ;
input   di ;
input   sr ;
input   en ;
input   clk ;

wire clk_in;
wire reset;
wire reg_enable;
reg qx;

initial begin
    qx = init;
end

assign reg_enable    = (always_en == 1'b1) ? 1'b1 : (en_inv == 1'b0) ? en : ~en;
assign clk_in     = (clk_inv == 1'b0) ? clk : ~clk;
assign reset    = (no_sr == 1'b1) ? 1'b0 : ((sr_inv == 1'b0) ? sr : ~sr);

if(latch_mode == 1'b1) begin
    always @ (*) begin
        if(reset)  
            qx <= sr_value;
        else if(reg_enable & clk_in)  
            qx <= di;
    end
end
else begin
    if(sync_mode == 1'b0) begin
        always @(posedge clk_in or posedge reset) begin
            if(reset)
                qx <= sr_value;
            else 
                if (reg_enable) begin
                    qx <= di;
                end
        end
    end else begin
        always @(posedge clk_in) begin
            if(reset)
                qx <= sr_value;
            else 
                if (reg_enable) begin
                    qx <= di;
                end
        end
    end
end

endmodule


module VCC (Y);
    output Y;

    assign Y = 1;
endmodule


module LRAM32X2SP(
input clk, 
input we, 
input [4:0] addr, 
input [1:0] din,  
output [1:0] dout 
); 

`ifdef  SIMULATION
    reg [63:0] config_data = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg    [1:0] ram [31:0];

integer count;

initial begin
    # 1;
    for(count = 0; count <32; count = count + 1) begin
        ram[count] = {config_data[count + 32], config_data[count]};
    end
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addr] <= din;
end

assign dout = ram[addr];

endmodule

module LRAM32X2QP(
    input clk, 
    input we, 
    input [4:0] addra, 
    input [4:0] addrb, 
    input [4:0] addrc, 
    input [4:0] addrd, 
    input[1:0] din, 
    output [1:0] douta, 
    output [1:0] doutb, 
    output [1:0] doutc, 
    output [1:0] doutd 
);

`ifdef  SIMULATION
    reg [63:0] config_data = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg    [1:0] ram [31:0];

integer count, baseaddr;

initial begin
    # 1;
    for(count = 0; count <32; count = count + 1) begin
        ram[count] = {config_data[count + 32], config_data[count]};
    end
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addra] <= din;
end

assign douta = ram[addra];
assign doutb = ram[addrb];
assign doutc = ram[addrc];
assign doutd = ram[addrd];

endmodule

module LRAM32M(
    input clk, 
    input we, 
    input [4:0] addra, 
    input [4:0] addrb, 
    input [4:0] addrc, 
    input [4:0] addrd, 
    input [1:0] dina, 
    input [1:0] dinb, 
    input [1:0] dinc, 
    input [1:0] dind, 
    output [1:0] douta, 
    output [1:0] doutb, 
    output [1:0] doutc, 
    output [1:0] doutd 
);

`ifdef  SIMULATION
    reg [63:0] config_data_a = 64'h0000_0000_0000_0000;
    reg [63:0] config_data_b = 64'h0000_0000_0000_0000;
    reg [63:0] config_data_c = 64'h0000_0000_0000_0000;
    reg [63:0] config_data_d = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data_a = 64'h0000_0000_0000_0000;    
    parameter config_data_b = 64'h0000_0000_0000_0000;    
    parameter config_data_c = 64'h0000_0000_0000_0000;    
    parameter config_data_d = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg    [1:0] rama [31:0];
reg    [1:0] ramb [31:0];
reg    [1:0] ramc [31:0];
reg    [1:0] ramd [31:0];

integer counta;
integer countb;
integer countc;
integer countd;

initial begin
    # 1;
    for(counta = 0; counta <32; counta = counta + 1) begin
        rama[counta] = {config_data_a[counta + 32], config_data_a[counta]};
    end
    for(countb = 0; countb <32; countb = countb + 1) begin
        ramb[countb] = {config_data_b[countb + 32], config_data_b[countb]};
    end
    for(countc = 0; countc <32; countc = countc + 1) begin
        ramc[countc] = {config_data_c[countc + 32], config_data_c[countc]};
    end
    for(countd = 0; countd <32; countd = countd + 1) begin
        ramd[countd] = {config_data_d[countd + 32], config_data_d[countd]};
    end
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we) begin
    rama[addra] <= dina;
    ramb[addra] <= dinb;
    ramc[addra] <= dinc;
    ramd[addra] <= dind;
end
end

assign douta = rama[addra];
assign doutb = ramb[addrb];
assign doutc = ramc[addrc];
assign doutd = ramd[addrd];

endmodule

module LRAM64X1SP(
input clk, 
input we, 
input [5:0] addr, 
input  din,  
output  dout 
); 

`ifdef  SIMULATION
    reg [63:0] config_data = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [63:0] ram;


initial begin
    # 1;
    ram = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addr] <= din;
end

assign dout = ram[addr];

endmodule

module LRAM64X1DP(
input clk, 
input we, 
input [5:0] addra, 
input [5:0] addrb, 
input  din,  
output  douta,
output  doutb 
); 

`ifdef  SIMULATION
    reg [63:0] config_data = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [63:0] ram;


initial begin
    # 1;
    ram = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addra] <= din;
end

assign douta = ram[addra];
assign doutb = ram[addrb];

endmodule

module LRAM64X1QP(
input clk, 
input we, 
input [5:0] addra, 
input [5:0] addrb, 
input [5:0] addrc, 
input [5:0] addrd, 
input  din,  
output  douta,
output  doutb,
output  doutc,
output  doutd 
); 

`ifdef  SIMULATION
    reg [63:0] config_data = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [63:0] ram;


initial begin
    # 1;
    ram = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addra] <= din;
end

assign douta = ram[addra];
assign doutb = ram[addrb];
assign doutc = ram[addrc];
assign doutd = ram[addrd];

endmodule

module LRAM64M(
input clk, 
input we, 
input [5:0] addra, 
input [5:0] addrb, 
input [5:0] addrc, 
input [5:0] addrd, 
input  dina,  
input  dinb,  
input  dinc,  
input  dind,  
output  douta,
output  doutb,
output  doutc,
output  doutd 
); 

`ifdef  SIMULATION
    reg [63:0] config_data_a = 64'h0000_0000_0000_0000;
    reg [63:0] config_data_b = 64'h0000_0000_0000_0000;
    reg [63:0] config_data_c = 64'h0000_0000_0000_0000;
    reg [63:0] config_data_d = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data_a = 64'h0000_0000_0000_0000;    
    parameter config_data_b = 64'h0000_0000_0000_0000;    
    parameter config_data_c = 64'h0000_0000_0000_0000;    
    parameter config_data_d = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [63:0] rama;
reg [63:0] ramb;
reg [63:0] ramc;
reg [63:0] ramd;


initial begin
    # 1;
    rama = config_data_a;
    ramb = config_data_b;
    ramc = config_data_c;
    ramd = config_data_d;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we) begin
    rama[addra] <= dina;
    ramb[addra] <= dinb;
    ramc[addra] <= dinc;
    ramd[addra] <= dind;
end
end

assign douta = rama[addra];
assign doutb = ramb[addrb];
assign doutc = ramc[addrc];
assign doutd = ramd[addrd];

endmodule

module LRAM128X1SP(
input clk, 
input we, 
input [6:0] addr, 
input  din,  
output  dout 
); 

`ifdef  SIMULATION
    reg [127:0] config_data = 128'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 128'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [127:0] ram;


initial begin
    # 1;
    ram = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addr] <= din;
end

assign dout = ram[addr];

endmodule

module LRAM128X2SP(
input clk, 
input we, 
input [6:0] addr, 
input  [1:0] din,  
output  [1:0] dout 
); 

`ifdef  SIMULATION
    reg [127:0] config_data_0 = 128'h0000_0000_0000_0000_0000_0000_0000_0000;
    reg [127:0] config_data_1 = 128'h0000_0000_0000_0000_0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data_0 = 128'h0000_0000_0000_0000_0000_0000_0000_0000;    
    parameter config_data_1 = 128'h0000_0000_0000_0000_0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [127:0] raml;
reg [127:0] ramh;


initial begin
    # 1;
    raml = config_data_0;
    ramh = config_data_1;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we) begin
    raml[addr] <= din[0];
    ramh[addr] <= din[1];
end
end

assign dout[0] = raml[addr];
assign dout[1] = ramh[addr];

endmodule

module LRAM128X1DP(
input clk, 
input we, 
input [6:0] addra, 
input [6:0] addrb, 
input  din,  
output  douta,
output  doutb 
); 

`ifdef  SIMULATION
    reg [127:0] config_data = 128'h0000_0000_0000_0000_0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 128'h0000_0000_0000_0000_0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [127:0] ram;


initial begin
    # 1;
    ram = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
if (we)
    ram[addra] <= din;
end

assign douta = ram[addra];
assign doutb = ram[addrb];

endmodule

module LRAM256X1SP(
input clk, 
input we, 
input [7:0] addr, 
input  din,  
output  dout 
); 

`ifdef  SIMULATION
    reg [255:0] config_data = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    parameter clk_inv = 1'b0;
`endif

reg [255:0] ram;

initial begin
    # 1;
    ram = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;


always @(posedge clk_in) begin
if (we)
    ram[addr] <= din;
end

assign dout = ram[addr];

endmodule

module SR16X2(
input [1:0] din,
input [3:0] addr,
input ce,
input clk,
output [1:0] dout
);


`ifdef  SIMULATION
    reg [15:0] config_data_h = 16'h0000;
    reg [15:0] config_data_l = 16'h0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data_h = 16'h0000;    
    parameter config_data_l = 16'h0000;    
    parameter clk_inv = 1'b0;
`endif

reg [15:0] SR_h;
reg [15:0] SR_l;

initial begin
    # 1;
    SR_h = config_data_h;
    SR_l = config_data_l;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
    if(ce) begin
        SR_h<= {SR_h[14:0], din[1]};
        SR_l<= {SR_l[14:0], din[0]};
    end
end

assign dout[1] = SR_h[addr];
assign dout[0] = SR_l[addr];

endmodule


module SR32X1(
input din,
input [4:0] addr,
input ce,
input clk,
output dout,
output shiftout
);


`ifdef  SIMULATION
    reg [31:0] config_data = 32'h0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 32'h0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [31:0] SR;

initial begin
    # 1;
    SR = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
    if(ce) begin
        SR<= {SR[30:0], din};
    end
end

assign shiftout = SR[31];
assign dout = SR[addr];

endmodule


module SR64X1(
input din,
input [5:0] addr,
input ce,
input clk,
output dout,
output shiftout
);


`ifdef  SIMULATION
    reg [63:0] config_data = 64'h0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 64'h0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [63:0] SR;

initial begin
    # 1;
    SR = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
    if(ce) begin
        SR<= {SR[62:0], din};
    end
end

assign shiftout = SR[63];
assign dout = SR[addr];

endmodule


module SR128X1(
input din,
input [6:0] addr,
input ce,
input clk,
output dout,
output shiftout
);


`ifdef  SIMULATION
    reg [127:0] config_data = 128'h0000_0000_0000_0000_0000_0000_0000_0000;
    reg clk_inv = 1'b0;
`else
    parameter config_data = 128'h0000_0000_0000_0000_0000_0000_0000_0000;    
    parameter clk_inv = 1'b0;
`endif

reg [127:0] SR;

initial begin
    # 1;
    SR = config_data;
end

wire clk_in = (clk_inv == 1'b0) ? clk : ~clk;

always @(posedge clk_in) begin
    if(ce) begin
        SR<= {SR[126:0], din};
    end
end

assign shiftout = SR[127];
assign dout = SR[addr];

endmodule

module GBUF(in, out);
    input in;
    output out;
    
    buf (out, in);
    
endmodule

module RBUF(in, out);
    input in;
    output out;
    
    buf (out, in);
    
endmodule

module DBUF(in, out);
    input in;
    output out;
    
    buf (out, in);
    
endmodule

module GBUF_GATE (
    clk,
    en,
    clk_out
);

    input clk;
    input en;
    output clk_out;
    
    reg en_latch;
    always @(*) begin
        if (clk == 0)
            en_latch <= en;
    end

    assign clk_out = clk & en_latch;

endmodule

module RBUF_GATE (
    clk,
    en,
    clk_out
);

    input clk;
    input en;
    output clk_out;
    
    reg en_latch;
    always @(*) begin
        if (clk == 0)
            en_latch <= en;
    end

    assign clk_out = clk & en_latch;

endmodule

module DBUF_GATE (
    clk,
    en,
    clk_out
);

    input clk;
    input en;
    output clk_out;

    reg en_latch;
    always @(*) begin
        if (clk == 0)
            en_latch <= en;
    end

    assign clk_out = clk & en_latch;

endmodule

module DELAY_BUF (
    in, 
    out
);

    input in ;
    output out ;
   
    buf (out, in);

endmodule

module MULT_18X18(R, A, B);
    
input signed     [17:0] A;
input signed     [17:0] B;
output signed   [35:0] R;

//Function    // multiplier
    assign R= A * B;

endmodule

module UNSIGNED_18X18(A, B, R);

  input [17:0] A;
  input [17:0] B;
  output [35:0] R;

//Function    // multiplier
    assign R= A * B;

endmodule

module MULT_35X18(R, A, B);
     
input signed     [34:0] A;
input signed     [17:0] B;
output signed    [52:0] R;

//Function    // multiplier
    assign R= A * B;

endmodule

module MULT_35X35(R, A, B);
    
input signed     [34:0] A;
input signed     [34:0] B;
output signed    [69:0] R;

//Function    // multiplier
    assign R= A * B;

endmodule

module MULT_69X18(A, B, R);

input signed     [68:0] A;
input signed     [17:0] B;
output signed    [86:0] R;

//Function    // multiplier
    assign R= A * B;

endmodule

module MULT_69X69(A, B, R);

input signed     [68:0] A;
input signed     [68:0] B;
output signed    [137:0] R;

//Function    // multiplier
    assign R= A * B;

endmodule

module EMB5K (doa, dob, dopa, dopb, 
             addra, addrb, clka, clkb, dia, dib, dipa, dipb, cea, ceb, regcea, regceb, 
             regsra, regsrb, wea, web);

    output [15:0] doa;
    output [7:0] dob;
    output [1:0] dopa;
    output [0:0] dopb;
    
    input cea, clka, regcea;
    input ceb, clkb, regceb;
    input regsra, regsrb;
    input [11:0] addra;
    input [11:0] addrb;
    input [15:0] dia;
    input [15:0] dib;
    input [1:0] dipa;
    input [1:0] dipb;
    input [0:0] wea;
    input [0:0] web;

    parameter outreg_a = 1'b0;
    parameter outreg_b = 1'b0;
    parameter writemode_a = "write_first";
    parameter writemode_b = "write_first";
    parameter width_a = 1;//0;
    parameter width_b = 0;
    parameter clka_inv = 1'b0;
    parameter clkb_inv = 1'b0;
    parameter rammode = "sdp";
    
    parameter init_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

    parameter init_file = "none";     

    localparam [3:0] modea_sel = (width_a == 1) ? 4'b1111 : 
                           (width_a == 2) ? 4'b1110 :
                           (width_a == 4) ? 4'b1100 :
                           (width_a == 9) ? 4'b1000 :
                           (width_a == 18) ? 4'b0000 : 4'bxxxx;
                           
    localparam [3:0] modeb_sel = (width_b == 1) ? 4'b1111 : 
                           (width_b == 2) ? 4'b1110 :
                           (width_b == 4) ? 4'b1100 :
                           (width_b == 9) ? 4'b1000 :
                           (width_b == 18) ? 4'b0000 : 4'bxxxx;

    localparam [1:0] modea_wr = (writemode_a == "write_first") ? 2'b01 :
                          (writemode_a == "no_change") ? 2'b00 :
                          (writemode_a == "read_first") ? 2'b11 : 2'bxx;
                          
    localparam [1:0] modeb_wr = (writemode_b == "write_first") ? 2'b01 :
                          (writemode_b == "no_change") ? 2'b00 :
                          (writemode_b == "read_first") ? 2'b11 : 2'bxx;                          
    
    wire [17:0] dataina = (width_a == 18) ? {dipa, dia} : 
                          (width_a == 9) ? {dipa[0], dipa[0], dia[7:0], dia[7:0]} :
                          (width_a == 4) ? {1'bx, 1'bx, {4{dia[3:0]}}} :
                          (width_a == 2) ? {1'bx, 1'bx, {8{dia[1:0]}}} :
                          (width_a == 1) ? {1'bx, 1'bx, {16{dia[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;
                          
    wire [17:0] datainb = (width_b == 18) ? {dipb, dib} : 
                          (width_b == 9) ? {dipb[0], dipb[0], dib[7:0], dib[7:0]} :
                          (width_b == 4) ? {1'bx, 1'bx, {4{dib[3:0]}}} :
                          (width_b == 2) ? {1'bx, 1'bx, {8{dib[1:0]}}} :
                          (width_b == 1) ? {1'bx, 1'bx, {16{dib[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;
  
    wire [17:0] dataout;
    
    wire [1:0] regen = (rammode == "tdp") ? {regceb, regcea} : {regcea, regcea};
    
    integer i;
    
    assign dopb = dataout[17];
    assign dopa[1] = dataout[17];
    assign dopa[0] = (width_a == 18) ? dataout[16] : dataout[8];
    assign dob = dataout[16:9];
    assign doa = dataout[15:0];
    // address translation
               
    //sp mode
    localparam sp_addr_lbit = (width_a == 1) ? 0 : (width_a == 2) ? 1 : 
                              (width_a == 4) ? 2 : (width_a == 9) ? 3 : 
                              (width_a == 18) ? 4 : 0; 
    //sdp mode
    localparam sdp_raddr_lbit = (width_a == 1) ? 0 : (width_a == 2) ? 1 : 
                                (width_a == 4) ? 2 : (width_a == 9) ? 3 : 
                                (width_a == 18) ? 4: 0;                 
    localparam sdp_waddr_lbit = (width_b == 1) ? 0 : (width_b == 2) ? 1 : 
                                (width_b == 4) ? 2 : (width_b == 9) ? 3 : 
                                (width_b == 18) ? 4 : 0; 
    //tdp mode
    localparam tdp_addra_lbit = (width_a == 1) ? 0 : (width_a == 2) ? 1 : 
                                (width_a == 4) ? 2 : (width_a == 9) ? 3 : 0;                   
    localparam tdp_addrb_lbit = (width_b == 1) ? 0 : (width_b == 2) ? 1 : 
                                (width_b == 4) ? 2 : (width_b == 9) ? 3 : 0;

    localparam addra_lbit = (rammode == "sp")  ? sp_addr_lbit :
                            (rammode == "sdp") ? sdp_raddr_lbit :
                            (rammode == "tdp") ? tdp_addra_lbit : 0;
    localparam addrb_lbit = (rammode == "sp")  ? sp_addr_lbit :
                            (rammode == "sdp") ? sdp_waddr_lbit :
                            (rammode == "tdp") ? tdp_addrb_lbit : 0;
    //translation
    wire [11:0] addra_input;
    wire [11:0] addrb_input;
    
    localparam  addr_width_a = (width_a == 1) ? 12 : (width_a == 2) ? 11 :
                               (width_a == 4) ? 10 : (width_a == 8) ? 9 :
                               (width_a == 9) ? 9 : (width_a == 16) ? 8 :
                               (width_a == 18) ? 8 : 0;
    localparam  addr_width_b = (width_b == 1) ? 12 : (width_b == 2) ? 11 :
                               (width_b == 4) ? 10 : (width_b == 8) ? 9 :
                               (width_b == 9) ? 9 : (width_b == 16) ? 8 :
                               (width_b == 18) ? 8 : 1;//sp mode not use port b default 1 for addrb_input[addrb_lbit + addr_width_b - 1 : addrb_lbit] = addrb; when with_b=0
                               
    assign addra_input[addra_lbit + addr_width_a - 1 : addra_lbit] = addra;    
    if (addra_lbit > 0)
        assign addra_input[addra_lbit - 1 : 0] = 0;
    if (addra_lbit + addr_width_a < 12)
        assign addra_input[11 : addra_lbit + addr_width_a] = 0;
        
    assign addrb_input[addrb_lbit + addr_width_b - 1 : addrb_lbit] = addrb;
    if (addrb_lbit > 0)
        assign addrb_input[addrb_lbit - 1 : 0] = 0;
    if (addrb_lbit + addr_width_b < 12)
        assign addrb_input[11 : addrb_lbit + addr_width_b] = 0; 
 
    
BRAM18KV1 # (
    .DEPTH_EXT_MODE23       (1'b0),
    .DEPTH_EXT_MODE01       (1'b0),
    .ECC_DEC_EN             (1'b0),
    .ECC_ENC_EN             (1'b0),    

    .EMB5K_4_MODEA_SEL      (),
    .EMB5K_4_MODEB_SEL      (),
    .EMB5K_4_PORTA_BYPASS   (),
    .EMB5K_4_PORTA_CE       (),
    .EMB5K_4_PORTA_REG_OUT  (),
    .EMB5K_4_PORTA_WR_MODE  (),
    .EMB5K_4_PORTA_CKINV    (),
    .EMB5K_4_PORTB_BYPASS   (),
    .EMB5K_4_PORTB_CE       (),
    .EMB5K_4_PORTB_REG_OUT  (),
    .EMB5K_4_PORTB_WR_MODE  (),
    .EMB5K_4_PORTB_CKINV    (),
    
    .EMB5K_3_MODEA_SEL      (),
    .EMB5K_3_MODEB_SEL      (),
    .EMB5K_3_PORTA_BYPASS   (),
    .EMB5K_3_PORTA_CE       (),
    .EMB5K_3_PORTA_REG_OUT  (),
    .EMB5K_3_PORTA_WR_MODE  (),
    .EMB5K_3_PORTA_CKINV    (),
    .EMB5K_3_PORTB_BYPASS   (),
    .EMB5K_3_PORTB_CE       (),
    .EMB5K_3_PORTB_REG_OUT  (),
    .EMB5K_3_PORTB_WR_MODE  (),
    .EMB5K_3_PORTB_CKINV    (),
    
    .EMB5K_2_MODEA_SEL      (),
    .EMB5K_2_MODEB_SEL      (),
    .EMB5K_2_PORTA_BYPASS   (),
    .EMB5K_2_PORTA_CE       (),
    .EMB5K_2_PORTA_REG_OUT  (),
    .EMB5K_2_PORTA_WR_MODE  (),
    .EMB5K_2_PORTA_CKINV    (),
    .EMB5K_2_PORTB_BYPASS   (),
    .EMB5K_2_PORTB_CE       (),
    .EMB5K_2_PORTB_REG_OUT  (),
    .EMB5K_2_PORTB_WR_MODE  (),
    .EMB5K_2_PORTB_CKINV    (),
    
    .EMB5K_1_MODEA_SEL      (modea_sel),
    .EMB5K_1_MODEB_SEL      (modeb_sel),
    .EMB5K_1_PORTA_BYPASS   (1'b0),
    .EMB5K_1_PORTA_CE       (1'b1),
    .EMB5K_1_PORTA_REG_OUT  (outreg_a),
    .EMB5K_1_PORTA_WR_MODE  (modea_wr),
    .EMB5K_1_PORTA_CKINV    (clka_inv),
    .EMB5K_1_PORTB_BYPASS   (1'b0),
    .EMB5K_1_PORTB_CE       (1'b1),
    .EMB5K_1_PORTB_REG_OUT  (outreg_b),
    .EMB5K_1_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_1_PORTB_CKINV    (clkb_inv),
    
    .EXT_18K                (1'b0),
    .FIFO_EN                (1'b0),
    .PORTA_PROG             (8'b11110000),
    .PORTB_PROG             (8'b00001111),
    .WIDTH_EXT_MODE23       (1'b0),
    .WIDTH_EXT_MODE01       (1'b0)
)

u0_emb18k_core (
    .a_addr_ext             (2'b00),
    .b_addr_ext             (2'b00),
    
    .c1r4_aa                (),
    .c1r4_ab                (),
    .c1r4_cea               (),
    .c1r4_ceb               (),
    .c1r4_clka              (),
    .c1r4_clkb              (),
    .c1r4_da                (),
    .c1r4_db                (),
    .c1r4_rstna             (),
    .c1r4_rstnb             (),
    .c1r4_wea               (),
    .c1r4_web               (),
    .c1r4_user_ena          (),
    .c1r4_user_enb          (),
    
    .c1r3_aa                (),
    .c1r3_ab                (),
    .c1r3_cea               (),
    .c1r3_ceb               (),
    .c1r3_clka              (),
    .c1r3_clkb              (),
    .c1r3_da                (),
    .c1r3_db                (),
    .c1r3_rstna             (),
    .c1r3_rstnb             (),
    .c1r3_wea               (),
    .c1r3_web               (),
    .c1r3_user_ena          (),
    .c1r3_user_enb          (),
    
    .c1r2_aa                (),
    .c1r2_ab                (),
    .c1r2_cea               (),
    .c1r2_ceb               (),
    .c1r2_clka              (),
    .c1r2_clkb              (),
    .c1r2_da                (),
    .c1r2_db                (),
    .c1r2_rstna             (),
    .c1r2_rstnb             (),
    .c1r2_wea               (),
    .c1r2_web               (),
    .c1r2_user_ena          (),
    .c1r2_user_enb          (),    
    
    .c1r1_aa                (addra_input),
    .c1r1_ab                (addrb_input),
    .c1r1_cea               (cea),
    .c1r1_ceb               (ceb),
    .c1r1_clka              (clka),
    .c1r1_clkb              (clkb),
    .c1r1_da                (dataina),
    .c1r1_db                (datainb),
    .c1r1_rstna             (regsra),
    .c1r1_rstnb             (regsrb),
    .c1r1_wea               (wea[0]),
    .c1r1_web               (web[0]),
    .c1r1_user_ena          (regen[0]),
    .c1r1_user_enb          (regen[1]),
    
    .rd_mem_n               (1'b0),
    .rptr                   (14'b0),
    .wptr                   (14'b0),
    .wr_mem_n               (1'b0),
        
    .c1r4_q                 (),
    .c1r3_q                 (),
    .c1r2_q                 (),
    .c1r1_q                 (dataout),
    .eccindberr             (1'b0),
    .eccinsberr             (1'b0),
    .eccoutdberr            (),
    .eccoutsberr            (),
    .err_addr               () 
);

wire GSR;
glbsr inst( .GSR( GSR )) ;

initial
begin
    @(posedge GSR);
    for (i = 0; i < 16; i = i + 1)
    begin
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i    ] <= {initp_00[i*2+1   -:2 ], init_00[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+16 ] <= {initp_00[i*2+33  -:2 ], init_01[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+32 ] <= {initp_00[i*2+65  -:2 ], init_02[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+48 ] <= {initp_00[i*2+97  -:2 ], init_03[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+64 ] <= {initp_00[i*2+129 -:2 ], init_04[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+80 ] <= {initp_00[i*2+161 -:2 ], init_05[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+96 ] <= {initp_00[i*2+193 -:2 ], init_06[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+112] <= {initp_00[i*2+225 -:2 ], init_07[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+128] <= {initp_01[i*2+1   -:2 ], init_08[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+144] <= {initp_01[i*2+33  -:2 ], init_09[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+160] <= {initp_01[i*2+65  -:2 ], init_0a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+176] <= {initp_01[i*2+97  -:2 ], init_0b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+192] <= {initp_01[i*2+129 -:2 ], init_0c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+208] <= {initp_01[i*2+161 -:2 ], init_0d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+224] <= {initp_01[i*2+193 -:2 ], init_0e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+240] <= {initp_01[i*2+225 -:2 ], init_0f[i*16+15 -:16 ]};
    end
end
  
endmodule // EMB5K

// end of EMB5K 

module EMB9K (doa, dob, dopa, dopb, 
             addra, addrb, clka, clkb, dia, dib, dipa, dipb, cea, ceb, regcea, regceb, 
             regsra, regsrb, wea, web);

    output [31:0] doa;
    output [15:0] dob;
    output [3:0] dopa;
    output [1:0] dopb;
    
    input cea, clka, regcea;
    input ceb, clkb, regceb;
    input regsra, regsrb;
    input [12:0] addra;
    input [12:0] addrb;
    input [31:0] dia;
    input [31:0] dib;
    input [3:0] dipa;
    input [3:0] dipb;
    input [1:0] wea;
    input [1:0] web;

    parameter outreg_a = 0;
    parameter outreg_b = 0;
    parameter byte_write_enable = 0;
    parameter writemode_a = "write_first";
    parameter writemode_b = "write_first";
    parameter width_a = 1;//0;
    parameter width_b = 0;
    parameter extension_mode = "area";
    parameter clka_inv = 1'b0;
    parameter clkb_inv = 1'b0;
    
    parameter init_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;  

    parameter init_file = "none";
    parameter rammode = "sdp";  // "tdp", "sdp", "sp"
    parameter use_parity = 0;

    reg finish_error = 0;
    
    initial begin
    
        case (width_a)
            1: begin
                case (width_b)
                    0, 1, 2, 4, 9: ;
                    18 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9.", width_a);
                            finish_error = 1;
                        end
                    end
                    36 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                        end
                    end                
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            
            2, 4: begin
                case (width_b)
                    0, 1, 2, 4, 9, 18: ;
                    36 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            9: begin
                case (width_b)
                    0, 1, 2, 4, 9: ;
                    18 : begin
                        if (rammode == "tdp" && use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b is 9.", width_a);
                            finish_error = 1;
                        end
                    end
                    36 : begin
                        if (use_parity == 1) begin
                            if (rammode == "tdp") begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b is 9.", width_a);
                                finish_error = 1;
                            end
                            else begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 9, 18.", width_a);
                                finish_error = 1;
                            end
                        end
                        else if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b is 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            18: begin
                case (width_b)
                    1 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    0, 2, 4, 18: ;
                    9: begin
                        if (use_parity == 1 && rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b is 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    36: begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_a is 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            36: begin
                if (rammode == "tdp") begin
                    $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18.", width_a);
                    finish_error = 1;
                end
                else begin
                    case (width_b)
                    1: begin
                        $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_a are 2, 4, 9, 18, 36.", width_a);                   // end
                        finish_error = 1;
                    end
                    0, 2, 4, 18, 36: ;
                    9: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                    
                    default : begin
                        $display("Attribute Syntax Error : The attribute width_a on EMB9K instance %m is set to %d, Legal value for attribute width_b are 2, 4, 9, 18, 36.", width_a);
                        finish_error = 1;
                    end
                endcase
                end
            end
            default: begin
                if (rammode == "tdp") begin
                    $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18.", width_a);
                    finish_error = 1;
                end
                else begin
                    $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18, 36.", width_a);
                    finish_error = 1;
                end
            end
        endcase

        if (finish_error == 1)
            $finish;
    end // end initial
    
    parameter depth_extension = (width_a == 1) ? 1'b1 :
                                (width_a == 2) ?    ((width_b == 1) ? 1'b1 :
                                                    (width_b == 18 && rammode == "tdp") ? 1'b0 :
                                                    (width_b == 36) ? 1'b0 :
                                                    ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                (width_a == 4) ?     ((width_b == 1) ? 1'b1 :
                                                    (width_b == 18 && rammode == "tdp") ? 1'b0 :
                                                    (width_b == 36) ? 1'b0 :
                                                    ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                (width_a == 9) ?    ((width_b == 1) ? 1'b1 :
                                                    (width_b == 9 && use_parity == 1) ? 1'b1 :
                                                    (width_b == 18) ?   (rammode == "tdp") ? 1'b0 : 
                                                                        (use_parity == 1) ? 1'b1 :
                                                                        ((extension_mode == "area") ? 1'b0 : 1'b1) :
                                                    (width_b == 36) ? 1'b0 :
                                                    ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                (width_a == 18) ?   ((width_b == 1) ? 1'b1 :
                                                    (rammode == "tdp") ? 1'b0 :
                                                    (width_b == 9) ?     (use_parity == 1) ? 1'b1 :
                                                                        ((extension_mode == "area") ? 1'b0 : 1'b1) :
                                                    (width_b == 18) ?   (byte_write_enable == 1) ? 1'b0 :
                                                                        ((extension_mode == "area") ? 1'b0 : 1'b1) :
                                                    (width_b == 36) ? 1'b0 :
                                                    ((extension_mode == "area") ? 1'b0 :
                                                     (byte_write_enable == 1) ? 1'b0 :1'b1)) :                                                 
                                (width_a == 36) ? 1'b0 :
                                (extension_mode == "area") ? 1'b0 : 1'b1;
                                
    parameter width_extension = (depth_extension == 1'b1) ? 1'b0 : 1'b1;
    
    parameter width_a_5k =  (width_a == 1) ? 1 : 
                            (width_a == 2) ? ((depth_extension == 1'b0) ? 1 : 2) :
                            (width_a == 4) ? ((depth_extension == 1'b0) ? 2 : 4) :
                            (width_a == 9) ? ((depth_extension == 1'b0) ? 4 : 9) :
                            (width_a == 18) ? ((depth_extension == 1'b0) ? 9 : 18) :
                            (width_a == 36) ? 18 : 18;
                            
    parameter width_b_5k =  (width_b == 1) ? 1 : 
                            (width_b == 2) ? ((depth_extension == 1'b0) ? 1 : 2) :
                            (width_b == 4) ? ((depth_extension == 1'b0) ? 2 : 4) :
                            (width_b == 9) ? ((depth_extension == 1'b0) ? 4 : 9) :
                            (width_b == 18) ? ((depth_extension == 1'b0) ? 9 : 18) :
                            (width_b == 36) ? 18 : 18;

    localparam [3:0] modea_sel = (width_a_5k == 1) ? 4'b1111 : 
                           (width_a_5k == 2) ? 4'b1110 :
                           (width_a_5k == 4) ? 4'b1100 :
                           (width_a_5k == 9) ? 4'b1000 :
                           (width_a_5k == 18) ? 4'b0000 : 4'b0000;
    localparam [3:0] modeb_sel = (width_b_5k == 1) ? 4'b1111 : 
                           (width_b_5k == 2) ? 4'b1110 :
                           (width_b_5k == 4) ? 4'b1100 :
                           (width_b_5k == 9) ? 4'b1000 :
                           (width_b_5k == 18) ? 4'b0000 : 4'b0000;
                           
    localparam [1:0] modea_wr =   (writemode_a == "write_first") ? 2'b01 :
                            (writemode_a == "no_change") ? 2'b00 :
                            (writemode_a == "read_first") ? 2'b11 : 2'b11;
                          
    localparam [1:0] modeb_wr =   (writemode_b == "write_first") ? 2'b01 :
                            (writemode_b == "no_change") ? 2'b00 :
                            (writemode_b == "read_first") ? 2'b11 : 2'b11;

     wire [17:0] dataina_bnk1 = (width_a_5k == 18) ? ((depth_extension == 1'b1) ?  {dipa[1:0], dia[15:0]}:
                                                      (width_a_5k <= width_b_5k) ? {dipa[1:0], dia[15:0]}:
                                                      (width_b_5k == 1) ? {dipa[2],dipa[0],dia[30], dia[28], dia[26], dia[24], dia[22], dia[20], dia[18], dia[16],dia[14], dia[12], dia[10], dia[8], dia[6], dia[4], dia[2], dia[0]}:
                                                      (width_b_5k == 2) ? {dipa[2],dipa[0],dia[29:28],dia[25:24],dia[21:20],dia[17:16],dia[13:12],dia[9:8],dia[5:4],dia[1:0]}:
                                                      (width_b_5k == 4) ? {dipa[2],dipa[0],dia[27:24],dia[19:16],dia[11:8],dia[3:0]}:
                                                      (width_b_5k == 9) ? {dipa[2],dipa[0], dia[23:16], dia[7:0]}:{dipa[1:0], dia[15:0]}) : 
                               (width_a_5k == 9) ? ((depth_extension == 1'b1) ?  {dipa[0], dipa[0], dia[7:0], dia[7:0]} :
                                                      (width_a_5k <= width_b_5k) ? {dipa[0], dipa[0], dia[7:0], dia[7:0]} :
                                                      (width_b_5k == 1) ? {dipa[0],dipa[0],dia[14], dia[12], dia[10], dia[8], dia[6], dia[4], dia[2], dia[0],dia[14], dia[12], dia[10], dia[8], dia[6], dia[4], dia[2], dia[0]}:
                                                      (width_b_5k == 2) ? {dipa[0],dipa[0],dia[13:12],dia[9:8],dia[5:4],dia[1:0],dia[13:12],dia[9:8],dia[5:4],dia[1:0]}:
                                                      (width_b_5k == 4) ? {dipa[0],dipa[0],dia[11:8],dia[3:0],dia[11:8],dia[3:0]}:{dipa[0], dipa[0], dia[7:0], dia[7:0]}) : 
                               (width_a_5k == 4) ? {1'bx, 1'bx, {4{dia[3:0]}}} :
                               (width_a_5k == 2) ? {1'bx, 1'bx, {8{dia[1:0]}}} :
                               (width_a_5k == 1) ? {1'bx, 1'bx, {16{dia[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;

    wire [17:0] dataina_bnk2 = (width_a_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[3:2], dia[31:16]}:
                                                      (width_b_5k == 1) ? {dipa[3],dipa[1],dia[31], dia[29], dia[27], dia[25], dia[23], dia[21], dia[19], dia[17],dia[15], dia[13], dia[11], dia[9], dia[7], dia[5], dia[3], dia[1]}:
                                                      (width_b_5k == 2) ? {dipa[3],dipa[1],dia[31:30],dia[27:26],dia[23:22],dia[19:18],dia[15:14],dia[11:10],dia[7:6],dia[3:2]}:
                                                      (width_b_5k == 4) ? {dipa[3],dipa[1],dia[31:28],dia[23:20],dia[15:12],dia[7:4]}:
                                                      (width_b_5k == 9) ? {dipa[3],dipa[1], dia[31:24], dia[15:8]}:{dipa[3:2], dia[31:16]}) : 
                               (width_a_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[1], dipa[1], dia[15:8], dia[15:8]} :
                                                      (width_b_5k == 1) ? {dipa[1],dipa[1],dia[15], dia[13], dia[11], dia[9], dia[7], dia[5], dia[3], dia[1],dia[15], dia[13], dia[11], dia[9], dia[7], dia[5], dia[3], dia[1]}:
                                                      (width_b_5k == 2) ? {dipa[1],dipa[1],dia[15:14],dia[11:10],dia[7:6],dia[3:2],dia[15:14],dia[11:10],dia[7:6],dia[3:2]}:
                                                      (width_b_5k == 4) ? {dipa[1],dipa[1],dia[15:12],dia[7:4],dia[15:12],dia[7:4]}:{dipa[1], dipa[1], dia[15:8], dia[15:8]}) :
                               (width_a_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{dia[7:4]}}}) :
                               (width_a_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dia[3:2]}}}) :
                               (width_a_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dia[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;

                               
    wire [17:0] datainb_bnk1 = (width_b_5k == 18) ? ((depth_extension == 1'b1) ? {dipb[1:0], dib[15:0]}:
                                                      (width_b_5k <= width_a_5k) ? {dipb[1:0], dib[15:0]}:
                                                      (width_a_5k == 1) ? {dipb[2],dipb[0],dib[30], dib[28], dib[26], dib[24], dib[22], dib[20], dib[18], dib[16],dib[14], dib[12], dib[10], dib[8], dib[6], dib[4], dib[2], dib[0]}:
                                                      (width_a_5k == 2) ? {dipb[2],dipb[0],dib[29:28],dib[25:24],dib[21:20],dib[17:16],dib[13:12],dib[9:8],dib[5:4],dib[1:0]}:
                                                      (width_a_5k == 4) ? {dipb[2],dipb[0],dib[27:24],dib[19:16],dib[11:8],dib[3:0]}:
                                                      (width_a_5k == 9) ? {dipb[2],dipb[0], dib[23:16], dib[7:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (width_b_5k == 9) ? ((depth_extension == 1'b1) ? {dipb[0], dipb[0], dib[7:0], dib[7:0]} :
                                                      (width_b_5k <= width_a_5k) ? {dipb[0], dipb[0], dib[7:0], dib[7:0]} :
                                                      (width_a_5k == 1) ? {dipb[0],dipb[0],dib[14], dib[12], dib[10], dib[8], dib[6], dib[4], dib[2], dib[0],dib[14], dib[12], dib[10], dib[8], dib[6], dib[4], dib[2], dib[0]}:
                                                      (width_a_5k == 2) ? {dipb[0],dipb[0],dib[13:12],dib[9:8],dib[5:4],dib[1:0],dib[13:12],dib[9:8],dib[5:4],dib[1:0]}:
                                                      (width_a_5k == 4) ? {dipb[0],dipb[0],dib[11:8],dib[3:0],dib[11:8],dib[3:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (width_b_5k == 4) ? {1'bx, 1'bx, {4{dib[3:0]}}} :
                               (width_b_5k == 2) ? {1'bx, 1'bx, {8{dib[1:0]}}} :
                               (width_b_5k == 1) ? {1'bx, 1'bx, {16{dib[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;

    wire [17:0] datainb_bnk2 = (width_b_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[3:2], dib[31:16]}:
                                                      (width_a_5k == 1) ? {dipb[3],dipb[1],dib[31], dib[29], dib[27], dib[25], dib[23], dib[21], dib[19], dib[17],dib[15], dib[13], dib[11], dib[9], dib[7], dib[5], dib[3], dib[1]}:
                                                      (width_a_5k == 2) ? {dipb[3],dipb[1],dib[31:30],dib[27:26],dib[23:22],dib[19:18],dib[15:14],dib[11:10],dib[7:6],dib[3:2]}:
                                                      (width_a_5k == 4) ? {dipb[3],dipb[1],dib[31:28],dib[23:20],dib[15:12],dib[7:4]}:
                                                      (width_a_5k == 9) ? {dipb[3],dipb[1], dib[31:24], dib[15:8]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_b_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[1], dipb[1], dib[15:8], dib[15:8]} :
                                                      (width_a_5k == 1) ? {dipb[1],dipb[1],dib[15], dib[13], dib[11], dib[9], dib[7], dib[5], dib[3], dib[1],dib[15], dib[13], dib[11], dib[9], dib[7], dib[5], dib[3], dib[1]}:
                                                      (width_a_5k == 2) ? {dipb[1],dipb[1],dib[15:14],dib[11:10],dib[7:6],dib[3:2],dib[15:14],dib[11:10],dib[7:6],dib[3:2]}:
                                                      (width_a_5k == 4) ? {dipb[1],dipb[1],dib[15:12],dib[7:4],dib[15:12],dib[7:4]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{dib[7:4]}}}) :
                               (width_b_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dib[3:2]}}}) :
                               (width_b_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dib[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                            
    wire [17:0] dataout_bnk1;
    wire [17:0] dataout_bnk2;
    
    wire [1:0] regen = (rammode == "tdp") ? {regceb, regcea} : {regcea, regcea};
    
    integer i;

   // assign dopb = (depth_extension == 1'b1) ? {1'bx, dataout_bnk1[17]} : {dataout_bnk2[17], dataout_bnk1[17]};
                 

    //assign dopa[3] = (depth_extension == 1'b1) ? 1'bx:dataout_bnk2[17];
    //assign dopa[2] = (depth_extension == 1'b1) ? 1'bx:((width_b_5k >= width_a_5k) ? dataout_bnk2[16] :dataout_bnk1[17]);
    //assign dopa[1] = (depth_extension == 1'b1) ? dataout_bnk1[17] : ((width_b_5k >= width_a_5k) ? dataout_bnk1[17] :dataout_bnk2[16]);
    //assign dopa[0] = (width_a_5k == 18) ? dataout_bnk1[16] : dataout_bnk1[8];

    //assign dopa[3] = dataout_bnk2[17];
    //assign dopa[1] = dataout_bnk1[17];
    //assign dopa[2] = (depth_extension == 1'b1) ? 1'bx : ((width_a_5k == 18) ? dataout_bnk2[16] : dataout_bnk2[8]);
    //assign dopa[0] = (width_a_5k == 18) ? dataout_bnk1[16] : dataout_bnk1[8];

    assign dopa[3] = (depth_extension == 1'b1) ? 1'bx : dataout_bnk2[17];
    //assign dopa[1] = (depth_extension == 1'b1) ? dataout_bnk1[17] :((width_a_5k == width_b_5k) ? dataout_bnk1[17] :((width_a_5k == 18) ? dataout_bnk2[16] : dataout_bnk2[8]));
    assign dopa[1] = (depth_extension == 1'b1) ? dataout_bnk1[17] :((width_a_5k == 9) ? dataout_bnk2[8] :((width_a_5k == 18) ? ((width_b_5k == 18) ?dataout_bnk1[17]: dataout_bnk2[16]) : dataout_bnk2[8]));
    assign dopa[2] = (depth_extension == 1'b1) ? 1'bx : ((width_a_5k == width_b_5k) ? dataout_bnk2[16]:dataout_bnk1[17]);
    assign dopa[0] = (width_a_5k == 18) ? dataout_bnk1[16] : dataout_bnk1[8];

    //assign dob[7:0] = dataout_bnk1[16:9];
    //assign dob[15:8] = (depth_extension == 1'b1) ? 8'bxxxxxxxx : {dataout_bnk2[16:9]};

    assign doa = width_a_5k==1 ? {30'h0,dataout_bnk2[0],dataout_bnk1[0]} :
                 width_a_5k==2 ? {28'h0,dataout_bnk2[1:0],dataout_bnk1[1:0]} :
                 width_a_5k==4 ? {24'h0,dataout_bnk2[3:0],dataout_bnk1[3:0]} :
                 width_a_5k==9 ? ((depth_extension == 1'b1) ? {16'h0,dataout_bnk2[7:0],dataout_bnk1[7:0]} :
                                   (width_b_5k >= width_a_5k) ?{16'h0,dataout_bnk2[7:0],dataout_bnk1[7:0]} :                            
                                   (width_b_5k == 4) ? {dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (width_b_5k == 2) ? {dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (width_b_5k == 1) ? {dataout_bnk2[7],dataout_bnk1[7],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk2[0],dataout_bnk1[0]}:{dataout_bnk2[15:0],dataout_bnk1[15:0]  }) :
                 
                 width_a_5k==18 ? ((depth_extension == 1'b1) ? {dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (width_b_5k >= width_a_5k) ?{dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (width_b_5k == 9) ? {dataout_bnk2[15:8],dataout_bnk1[15:8],dataout_bnk2[7:0],dataout_bnk1[7:0]  }:
                                   (width_b_5k == 4) ? {dataout_bnk2[15:12],dataout_bnk1[15:12],dataout_bnk2[11:8],dataout_bnk1[11:8],dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (width_b_5k == 2) ? {dataout_bnk2[15:14],dataout_bnk1[15:14],dataout_bnk2[13:12],dataout_bnk1[13:12],dataout_bnk2[11:10],dataout_bnk1[11:10],dataout_bnk2[9:8],dataout_bnk1[9:8],dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (width_b_5k == 1) ? {dataout_bnk2[15],dataout_bnk1[15],dataout_bnk2[14],dataout_bnk1[14],dataout_bnk2[13],dataout_bnk1[13],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk2[9],dataout_bnk1[9],dataout_bnk2[8],dataout_bnk1[8],dataout_bnk2[7],dataout_bnk1[7],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk2[0],dataout_bnk1[0]}:{dataout_bnk2[15:0],dataout_bnk1[15:0]  }) :
                 32'hxxxx_xxxx;

    assign dopb = (depth_extension == 1'b1) ? {1'bx, dataout_bnk1[17]} : {dataout_bnk2[17], dataout_bnk1[17]};

    assign dob = width_b_5k==1 ? {14'h0,dataout_bnk2[9],dataout_bnk1[9]} :
                 width_b_5k==2 ? {12'h0,dataout_bnk2[10:9],dataout_bnk1[10:9]} :
                 width_b_5k==4 ? {8'h0,dataout_bnk2[12:9],dataout_bnk1[12:9]} :
                 width_b_5k==9 ? ((depth_extension == 1'b1) ? {dataout_bnk2[16:9],dataout_bnk1[16:9]} :
                                  (width_a_5k >= width_b_5k) ?{dataout_bnk2[16:9],dataout_bnk1[16:9]} :
                                  (width_a_5k == 4) ?{dataout_bnk2[16:13],dataout_bnk1[16:13],dataout_bnk2[12:9],dataout_bnk1[12:9]  }:
                                  (width_a_5k == 2) ?{dataout_bnk2[16:15],dataout_bnk1[16:15],dataout_bnk2[14:13],dataout_bnk1[14:13],dataout_bnk2[12:11],dataout_bnk1[12:11],dataout_bnk2[10:9],dataout_bnk1[10:9] }:
                                  (width_a_5k == 1) ?{dataout_bnk2[16],dataout_bnk1[16],dataout_bnk2[15],dataout_bnk1[15] ,dataout_bnk2[14],dataout_bnk1[14],dataout_bnk2[13],dataout_bnk1[13],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk2[9],dataout_bnk1[9] }:16'hxxxx):

                 16'hxxxx;  
                 
    // address translation
               
    //sp mode
    localparam sp_addr_lbit = (width_a == 1) ? 0 : (width_a == 2) ? 1 : 
                              (width_a == 4) ? 2 : (width_a == 9) ? 3 : 
                              (width_a == 18) ? ((byte_write_enable == 1) ? 3:4) : 
                              (width_a == 36) ? 4 : 0;
    //sdp mode
    localparam sdp_raddr_lbit = (width_a == 1) ? 0 : 
                                (width_a == 2) ? ((width_b == 36) ? 0:1) : 
                                (width_a == 4) ? ((width_b == 36) ? 1:2) : 
                                (width_a == 9) ? ((width_b == 36) ? 2:3) : 
                                (width_a == 18) ? ((byte_write_enable == 1) ? 3:
                                ((width_b == 36) ? 3:4)) : (width_a == 36) ? 4 : 0;
                       
    localparam sdp_waddr_lbit = (width_b == 1) ? 0 : 
                                (width_b == 2) ? ((width_a == 36) ? 0 : 1) : 
                                (width_b == 4) ? ((width_a == 36) ? 1 : 2) : 
                                (width_b == 9) ? ((width_a == 36) ? 2 : 3) : 
                                (width_b == 18) ? ((byte_write_enable == 1) ? 3:
                                ((width_a == 36) ? 3 : 4)) : (width_b == 36) ? 4 : 0; 
    //tdp mode
    localparam tdp_addra_lbit = (width_a == 1) ? 0 : 
                                (width_a == 2) ? ((width_b == 18) ? 0:1)  : 
                                (width_a == 4) ? ((width_b == 18) ? 1:2) : 
                                (width_a == 9) ? ((width_b == 18) ? 2:3) : 
                                (width_a == 18) ? 3: 0;
                       
    localparam tdp_addrb_lbit = (width_b == 1) ? 0 : 
                                (width_b == 2) ? ((width_a== 18) ? 0:1) : 
                                (width_b == 4) ? ((width_a== 18) ? 1:2) : 
                                (width_b == 9) ? ((width_a== 18) ? 2:3) : 
                                (width_b == 18) ? 3:  0;
                   

    localparam addra_lbit = (rammode == "sp")  ? sp_addr_lbit :
                            (rammode == "sdp") ? sdp_raddr_lbit :
                            (rammode == "tdp") ? tdp_addra_lbit : 0;
    localparam addrb_lbit = (rammode == "sp")  ? sp_addr_lbit :
                            (rammode == "sdp") ? sdp_waddr_lbit :
                            (rammode == "tdp") ? tdp_addrb_lbit : 0;
    //translation
    wire [12:0] addra_input;
    wire [12:0] addrb_input;
    
    localparam  addr_width_a = (width_a == 1) ? 13 : (width_a == 2) ? 12 :
                               (width_a == 4) ? 11 : (width_a == 8) ? 10 :
                               (width_a == 9) ? 10 : (width_a == 16) ? 9 :
                               (width_a == 18) ? 9 : (width_a == 32) ? 8 :
                               (width_a == 36) ? 8 : 0;
    localparam  addr_width_b = (width_b == 1) ? 13 : (width_b == 2) ? 12 :
                               (width_b == 4) ? 11 : (width_b == 8) ? 10 :
                               (width_b == 9) ? 10 : (width_b == 16) ? 9 :
                               (width_b == 18) ? 9 : (width_b == 32) ? 8 :
                               (width_b == 36) ? 8 : 1;//sp mode not use port b default 1 for addrb_input[addrb_lbit + addr_width_b - 1 : addrb_lbit] = addrb; when with_b=0
                               
    assign addra_input[addra_lbit + addr_width_a - 1 : addra_lbit] = addra;    
    if (addra_lbit > 0)
        assign addra_input[addra_lbit - 1 : 0] = 0;
    if (addra_lbit + addr_width_a < 13)
        assign addra_input[12 : addra_lbit + addr_width_a] = 0;
        
    assign addrb_input[addrb_lbit + addr_width_b - 1 : addrb_lbit] = addrb;
    if (addrb_lbit > 0)
        assign addrb_input[addrb_lbit - 1 : 0] = 0;
    if (addrb_lbit + addr_width_b < 13)
        assign addrb_input[12 : addrb_lbit + addr_width_b] = 0; 

                             
BRAM18KV1 # (
    .DEPTH_EXT_MODE23        (1'b0),
    .DEPTH_EXT_MODE01        (depth_extension),
    .ECC_DEC_EN                (1'b0),
    .ECC_ENC_EN                (1'b0),
    
    .EMB5K_4_MODEA_SEL      (),
    .EMB5K_4_MODEB_SEL      (),
    .EMB5K_4_PORTA_BYPASS   (),
    .EMB5K_4_PORTA_CE       (),
    .EMB5K_4_PORTA_REG_OUT  (),
    .EMB5K_4_PORTA_WR_MODE  (),
    .EMB5K_4_PORTA_CKINV    (),
    .EMB5K_4_PORTB_BYPASS   (),
    .EMB5K_4_PORTB_CE       (),
    .EMB5K_4_PORTB_REG_OUT  (),
    .EMB5K_4_PORTB_WR_MODE  (),
    .EMB5K_4_PORTB_CKINV    (),
    
    .EMB5K_3_MODEA_SEL      (),
    .EMB5K_3_MODEB_SEL      (),
    .EMB5K_3_PORTA_BYPASS   (),
    .EMB5K_3_PORTA_CE       (),
    .EMB5K_3_PORTA_REG_OUT  (),
    .EMB5K_3_PORTA_WR_MODE  (),
    .EMB5K_3_PORTA_CKINV    (),
    .EMB5K_3_PORTB_BYPASS   (),
    .EMB5K_3_PORTB_CE       (),
    .EMB5K_3_PORTB_REG_OUT  (),
    .EMB5K_3_PORTB_WR_MODE  (),
    .EMB5K_3_PORTB_CKINV    (),
    
    .EMB5K_2_MODEA_SEL      (modea_sel),
    .EMB5K_2_MODEB_SEL      (modeb_sel),
    .EMB5K_2_PORTA_BYPASS   (1'b0),
    .EMB5K_2_PORTA_CE       (1'b1),
    .EMB5K_2_PORTA_REG_OUT  (outreg_a),
    .EMB5K_2_PORTA_WR_MODE  (modea_wr),
    .EMB5K_2_PORTA_CKINV    (clka_inv),
    .EMB5K_2_PORTB_BYPASS   (1'b0),
    .EMB5K_2_PORTB_CE       (1'b1),
    .EMB5K_2_PORTB_REG_OUT  (outreg_b),
    .EMB5K_2_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_2_PORTB_CKINV    (clkb_inv),
    
    .EMB5K_1_MODEA_SEL      (modea_sel),
    .EMB5K_1_MODEB_SEL      (modeb_sel),
    .EMB5K_1_PORTA_BYPASS   (1'b0),
    .EMB5K_1_PORTA_CE       (1'b1),
    .EMB5K_1_PORTA_REG_OUT  (outreg_a),
    .EMB5K_1_PORTA_WR_MODE  (modea_wr),
    .EMB5K_1_PORTA_CKINV    (clka_inv),
    .EMB5K_1_PORTB_BYPASS   (1'b0),
    .EMB5K_1_PORTB_CE       (1'b1),
    .EMB5K_1_PORTB_REG_OUT  (outreg_b),
    .EMB5K_1_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_1_PORTB_CKINV    (clkb_inv),
    
    .EXT_18K                (1'b0),
    .FIFO_EN                (1'b0),
    .PORTA_PROG                (8'b11110000),
    .PORTB_PROG                (8'b00001111),
    .WIDTH_EXT_MODE23        (1'b0),
    .WIDTH_EXT_MODE01        (width_extension)
)

u0_emb18k_core (
    .a_addr_ext                ({1'b1, addra_input[12]}),
    .b_addr_ext                ({1'b1, addrb_input[12]}),
    
    .c1r4_aa                (),
    .c1r4_ab                (),
    .c1r4_cea                (),
    .c1r4_ceb                (),
    .c1r4_clka                (),
    .c1r4_clkb                (),
    .c1r4_da                (),
    .c1r4_db                (),
    .c1r4_rstna                (),
    .c1r4_rstnb                (),
    .c1r4_wea                (),
    .c1r4_web                (),
    .c1r4_user_ena          (),
    .c1r4_user_enb          (),    
    
    .c1r3_aa                (),
    .c1r3_ab                (),
    .c1r3_cea                (),
    .c1r3_ceb                (),
    .c1r3_clka                (),
    .c1r3_clkb                (),
    .c1r3_da                (),
    .c1r3_db                (),
    .c1r3_rstna                (),
    .c1r3_rstnb                (),
    .c1r3_wea                (),
    .c1r3_web                (),
    .c1r3_user_ena          (),
    .c1r3_user_enb          (),    
    
    .c1r2_aa                (addra_input[11:0]),
    .c1r2_ab                (addrb_input[11:0]),
    .c1r2_cea                (cea),
    .c1r2_ceb                (ceb),
    .c1r2_clka                (clka),
    .c1r2_clkb                (clkb),
    .c1r2_da                (dataina_bnk2),
    .c1r2_db                (datainb_bnk2),
    .c1r2_rstna                (regsra),
    .c1r2_rstnb                (regsrb),
    .c1r2_wea                (wea[1]),
    .c1r2_web                (web[1]),
    .c1r2_user_ena          (regen[0]),
    .c1r2_user_enb          (regen[1]),
    
    .c1r1_aa                (addra_input[11:0]),
    .c1r1_ab                (addrb_input[11:0]),
    .c1r1_cea                (cea),
    .c1r1_ceb                (ceb),
    .c1r1_clka                (clka),
    .c1r1_clkb                (clkb),
    .c1r1_da                (dataina_bnk1),
    .c1r1_db                (datainb_bnk1),
    .c1r1_rstna                (regsra),
    .c1r1_rstnb                (regsrb),
    .c1r1_wea                (wea[0]),
    .c1r1_web                (web[0]),
    .c1r1_user_ena          (regen[0]),
    .c1r1_user_enb          (regen[1]),    
    
    .rd_mem_n                (1'b0),
    .rptr                    (14'b0),
    .wptr                    (14'b0),
    .wr_mem_n                (1'b0),
        
    .c1r4_q                    (),
    .c1r3_q                    (),
    .c1r2_q                    (dataout_bnk2),
    .c1r1_q                    (dataout_bnk1),
    .eccindberr             (1'b0),
    .eccinsberr             (1'b0),
    .eccoutdberr            (),
    .eccoutsberr            (),
    .err_addr                () 
    );

wire GSR;
glbsr inst( .GSR( GSR )) ;

initial
begin
    @(posedge GSR);
    for (i = 0; i < 16; i = i + 1)
    begin
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i    ] <= {initp_00[i*2+1   -:2 ], init_00[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+16 ] <= {initp_00[i*2+33  -:2 ], init_01[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+32 ] <= {initp_00[i*2+65  -:2 ], init_02[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+48 ] <= {initp_00[i*2+97  -:2 ], init_03[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+64 ] <= {initp_00[i*2+129 -:2 ], init_04[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+80 ] <= {initp_00[i*2+161 -:2 ], init_05[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+96 ] <= {initp_00[i*2+193 -:2 ], init_06[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+112] <= {initp_00[i*2+225 -:2 ], init_07[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+128] <= {initp_01[i*2+1   -:2 ], init_08[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+144] <= {initp_01[i*2+33  -:2 ], init_09[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+160] <= {initp_01[i*2+65  -:2 ], init_0a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+176] <= {initp_01[i*2+97  -:2 ], init_0b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+192] <= {initp_01[i*2+129 -:2 ], init_0c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+208] <= {initp_01[i*2+161 -:2 ], init_0d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+224] <= {initp_01[i*2+193 -:2 ], init_0e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+240] <= {initp_01[i*2+225 -:2 ], init_0f[i*16+15 -:16 ]};
        
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i    ] <= {initp_02[i*2+1   -:2 ], init_10[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+16 ] <= {initp_02[i*2+33  -:2 ], init_11[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+32 ] <= {initp_02[i*2+65  -:2 ], init_12[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+48 ] <= {initp_02[i*2+97  -:2 ], init_13[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+64 ] <= {initp_02[i*2+129 -:2 ], init_14[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+80 ] <= {initp_02[i*2+161 -:2 ], init_15[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+96 ] <= {initp_02[i*2+193 -:2 ], init_16[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+112] <= {initp_02[i*2+225 -:2 ], init_17[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+128] <= {initp_03[i*2+1   -:2 ], init_18[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+144] <= {initp_03[i*2+33  -:2 ], init_19[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+160] <= {initp_03[i*2+65  -:2 ], init_1a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+176] <= {initp_03[i*2+97  -:2 ], init_1b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+192] <= {initp_03[i*2+129 -:2 ], init_1c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+208] <= {initp_03[i*2+161 -:2 ], init_1d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+224] <= {initp_03[i*2+193 -:2 ], init_1e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+240] <= {initp_03[i*2+225 -:2 ], init_1f[i*16+15 -:16 ]};
    end
end
    
endmodule // EMB9K

// end of EMB9K 

module EMB18K (doa, dob, dopa, dopb, 
             addra, addrb, clka, clkb, dia, dib, dipa, dipb, cea, ceb, regcea, regceb, 
             regsra, regsrb, wea, web, eccoutdberr, eccoutsberr, eccreadaddr, eccindberr, eccinsberr);

    output [63:0] doa;
    output [31:0] dob;
    output [7:0] dopa;
    output [3:0] dopb;
    output eccoutdberr, eccoutsberr;
    output [7:0] eccreadaddr;
    
    input cea, clka, regcea;
    input ceb, clkb, regceb;
    input regsra, regsrb;
    input [13:0] addra;
    input [13:0] addrb;
    input [63:0] dia;
    input [63:0] dib;
    input [7:0] dipa;
    input [7:0] dipb;
    input [3:0] wea;
    input [3:0] web;
    input eccindberr, eccinsberr;

    parameter eccreaden = 0;
    parameter eccwriteen = 0;
    parameter outreg_a = 0;
    parameter outreg_b = 0;
    parameter writemode_a = "write_first";  // "write_first", "read_first", "no_change"
    parameter writemode_b = "write_first";  // "write_first", "read_first", "no_change"
    parameter width_a = 1;//0;
    parameter width_b = 0;
    parameter clka_inv = 1'b0;
    parameter clkb_inv = 1'b0;
    parameter extension_mode = "power"; // "area", "power"
    parameter rammode = "sdp";  // "tdp", "sdp", "sp"
    parameter use_parity = 0;
    
    parameter init_file = "none";
    
    parameter init_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_1f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_2a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_2b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_2c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_2d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_2e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_2f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_3a = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_3b = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_3c = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_3d = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_3e = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_3f = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

    reg finish_error = 0;
    
    initial begin 
        case (width_a)
            1: begin
                case (width_b)
                    0, 1, 2, 4, 9: ;
                    18 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            
            2: begin
                case (width_b)
                    0, 1, 2, 4, 9, 18: ;
                    36 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            
            4: begin
                case (width_b)
                    0, 1, 2, 4, 9, 18, 36: ;
                    72 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36, 72.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            9: begin
                case (width_b)
                    0, 1, 2, 4, 9: ;
                    18 : begin
                        if (rammode == "tdp" && use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 9.", width_a);
                            finish_error = 1;
                        end
                    end
                    36 : begin
                        if (use_parity == 1) begin
                            if (rammode == "tdp") begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 9.", width_a);
                                finish_error = 1;
                            end
                            else begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 9, 18.", width_a);
                                finish_error = 1;
                            end
                        end                
                    end
                    
                    72 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36, 72.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            18: begin
                case (width_b)
                    1, 72 : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                    0, 2, 4, 18: ;
                    9, 36: begin
                        if (use_parity == 1 && rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 18.", width_a);
                            finish_error = 1;
                        end
                    end
                    72: begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 18.", width_a);
                            finish_error = 1;
                        end
                        else if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                    end
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 2, 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 1, 2, 4, 9, 18, 36, 72.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            36: begin
                case (width_b)
                    1, 2: begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                        //else begin
                        //    $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 4, 9, 18, 36, 72.", width_a);
                        //    finish_error = 1;
                        //end
                    end
                    0, 4, 36: ;
                    9: begin
                        if (use_parity == 1) begin
                            if (rammode == "tdp") begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 36.", width_a);
                                finish_error = 1;
                            end
                            else begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 18, 36, 72.", width_a);
                                finish_error = 1;
                            end
                        end
                    end
                    18: begin
                        if (use_parity == 1 && rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 36.", width_a);
                            finish_error = 1;
                        end                    
                    end
                    72: begin
                        if (rammode == "tdp") begin
                            if (use_parity == 1) begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b is 36.", width_a);
                                finish_error = 1;
                            end
                            else begin
                                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 4, 9, 18, 36.", width_a);
                                finish_error = 1;
                            end
                        end                     
                    end
                    
                    default : begin
                        if (rammode == "tdp") begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 4, 9, 18, 36.", width_a);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 2, 4, 9, 18, 36, 72.", width_a);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            72: begin
                if (rammode == "tdp") begin
                    $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18, 36.", width_a);
                    finish_error = 1;
                end
                else begin            
                    case (width_b)
                        1, 2 : begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 4, 9, 18, 36, 72.", width_a);
                            finish_error = 1;
                        end
                    
                        0, 4, 9, 18, 36, 72: ;
    
                        default : begin
                            $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_b are 4, 9, 18, 36, 72.", width_a);
                            finish_error = 1;
                        end
                    endcase
                end
            end
        default: begin
            if (rammode == "tdp") begin
                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18, 36.", width_a);
                finish_error = 1;
            end
            else begin
                $display("Attribute Syntax Error : The attribute width_a on EMB18K instance %m is set to %d, Legal value for attribute width_a are 1, 2, 4, 9, 18, 36, 72.", width_a);
                finish_error = 1;
            end
        end
        endcase
        
        if (finish_error == 1)
            $finish;
    end // end initial
    
    // parameter depth_extension_0 =   (width_a == 1) ? 1'b1 :
                                    // (width_a == 2) ? 1'b1 :
                                    // (width_a == 4) ?    ((width_b == 1) ? 1'b1 :
                                                        // (width_b == 2) ? 1'b1 :
                                                        // (width_b == 18 && rammode == "tdp") ? 1'b0 :
                                                        // (width_b == 36) ? 1'b0 :
                                                        // (width_b == 72) ? 1'b0 :
                                                        // ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                    // (width_a == 9) ?    ((width_b == 1) ? 1'b1 :
                                                        // (width_b == 2) ? 1'b1 :
                                                        // (width_b == 9 && use_parity == 1) ? 1'b1 :
                                                        // (width_b == 18) ?   (rammode == "tdp") ? 1'b1 : 
                                                                            // (use_parity == 1) ? 1'b1 : 
                                                                            // ((extension_mode == "area") ? 1'b0 : 1'b1) :
                                                        // (width_b == 36) ? 1'b0 :
                                                        // (width_b == 72) ? 1'b0 :
                                                        // ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                    // (width_a == 18) ?   ((width_b == 1) ? 1'b1 :
                                                        // (width_b == 2) ? 1'b1 :
                                                        // (width_b == 9 && rammode != "tdp" && use_parity == 1) ? 1'b1 :
                                                        // (width_b == 18 && use_parity == 1) ? 1'b1 :
                                                        // (width_b == 36) ? 1'b0 :
                                                        // (width_b == 72) ? 1'b0 :
                                                        // ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                    // (width_a == 36) ?   ((width_b == 2 && rammode != "tdp") ? 1'b1 : 1'b0) :
                                    // (width_a == 72) ?   1'b0 : 1'b0;
                                
    // parameter width_extension_0 =   (depth_extension == 1'b1) ? 1'b0 : 1'b1;
    
    // parameter depth_extension_1 =   (width_a == 1) ? 1'b1 :
                                    // (width_a == 2) ? ((width_b == 16 && rammode == "tdp") ? 1'b0 :
                                                     // (width_b == 32 && rammode != "tdp") ? 1'b0 :
                                                     // 1'b1) :
                                    // (width_a == 4) ? ((width_b == 1) ? 1'b1 :
                                                     // (width_b == 2) ? 1'b1 :
                                                     // (width_b == 18 && rammode == "tdp") ? 1'b0 :
                                                     // (width_b == 36) ? 1'b0 :
                                                     // (width_b == 72) ? 1'b0 :
                                                     // ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                    // (width_a == 9) ? ((width_b == 1) ? 1'b1 :
                                                     // (width_b == 2) ? 1'b1 :
                                                     // (width_b == 9 && use_parity == 1) ? 1'b1 :
                                                     // (width_b == 18) ? (rammode == "tdp") ? 1'b0 : 
                                                                       // (use_parity == 1) ? 1'b1 :
                                                                       // ((extension_mode == "area") ? 1'b0 : 1'b1) :
                                                     // (width_b == 36) ? 1'b0 :
                                                     // (width_b == 72) ? 1'b0 :
                                                     // ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                    // (width_a == 18) ? ((width_b == 2) ? ((rammode == "tdp") ? 1'b0 : 1'b1) :
                                                      // (width_b == 9 && rammode != "tdp" && use_parity == 1) ? 1'b1 :
                                                      // (width_b == 18 && use_parity == 1) ? ((rammode == "tdp") ? 1'b0 : 1'b1) :
                                                      // (width_b == 36) ? 1'b0 :
                                                      // (width_b == 72) ? 1'b0 :
                                                      // ((extension_mode == "area") ? 1'b0 : 1'b1)) :
                                    // (width_a == 36) ? 1'b0 :
                                    // (width_a == 72) ? 1'b0 : 1'b0;
                                    
    // parameter extension18k =    (depth_extension_1 == depth_extension_0) ? 1'b1 : 1'b0;
                                

    // parameter width_a_5k =  (width_a == 1) ? 1 : 
                            // (width_a == 2) ? ((depth_extension_1 == 1'b0) ? 1 : 2) :
                            // (width_a == 4) ? ((depth_extension_1 == 1'b0) ? ((depth_extension_0 == 1'b0) ? 1 : 2) : 4) :
                            // (width_a == 9) ? ((depth_extension_1 == 1'b0) ? ((depth_extension_0 == 1'b0) ? 2 : 4) : 9) :
                            // (width_a == 18) ? ((depth_extension_1 == 1'b0) ? ((depth_extension_0 == 1'b0) ? 4 : 9) : 18) :
                            // (width_a == 36) ? ((depth_extension_0 == 1'b0) ? 9 : 18) :
                            // (width_a == 72) ? 18 : 18;
                            
    // parameter width_b_5k =  (width_b == 1) ? 1 : 
                            // (width_b == 2) ? ((depth_extension_1 == 1'b0) ? 1 : 2) :
                            // (width_b == 4) ? ((depth_extension_1 == 1'b0) ? ((depth_extension_0 == 1'b0) ? 1 : 2) : 4) :
                            // (width_b == 9) ? ((depth_extension_1 == 1'b0) ? ((depth_extension_0 == 1'b0) ? 2 : 4) : 9) :
                            // (width_b == 18) ? ((depth_extension_1 == 1'b0) ? ((depth_extension_0 == 1'b0) ? 4 : 9) : 18) :
                            // (width_b == 36) ? ((depth_extension_0 == 1'b0) ? 9 : 18) :
                            // (width_b == 72) ? 18 : 18;                       
    parameter depth_extension =   (width_a == 1) ? 1'b1 :
                                  (width_a == 2) ? 1'b1 :
                                  (width_a == 4) ? ((width_b == 1) ? 1'b1 :
                                                    (width_b == 2) ? 1'b1 :
                                                    (width_b == 4) ? 1'b1 :
                                                    (width_b == 9) ? 1'b1 :
                                                    (width_b == 18 ) ? (rammode == "tdp") ? 1'b0 : 1'b1 :
                                                    (width_b == 36) ? 1'b0 :
                                                    (width_b == 72) ? 1'b0 :
                                                    1'b1) :
                                  (width_a == 9) ? ((width_b == 1) ? 1'b1 :
                                                    (width_b == 2) ? 1'b1 :
                                                    (width_b == 4) ? 1'b1 :
                                                    (width_b == 9) ? 1'b1 : 
                                                    (width_b == 18) ? (rammode == "tdp") ? 1'b0 : 1'b1 :
                                                    (width_b == 36) ? 1'b0 :
                                                    (width_b == 72) ? 1'b0 :
                                                    1'b1) :
                                  (width_a == 18) ? ((rammode == "tdp") ? 1'b0 : 
                                                     (width_b == 1) ? 1'b1 :
                                                     (width_b == 2) ? 1'b1 :
                                                     (width_b == 9) ? 1'b1 :
                                                     (width_b == 18) ? 1'b1 :
                                                     (width_b == 36) ? 1'b0 :
                                                     (width_b == 72) ? 1'b0 :
                                                     1'b1) :
                                  (width_a == 36) ? 1'b0 :
                                  (width_a == 72) ? 1'b0 : 1'b1;
                                
    parameter width_extension =   (depth_extension == 1'b1) ? 1'b0 : 1'b1;
    
                                    
    // parameter extension18k =    depth_extension || width_extension;
    parameter extension18k =    1'b1;
                                

    parameter width_a_5k =  (width_a == 1) ? 1 : 
                            (width_a == 2) ? 2 :
                            (width_a == 4) ? ((depth_extension == 1) ? 4 : 1) :
                            (width_a == 9) ? ((depth_extension == 1) ? 9 : 2) :
                            (width_a == 18) ? ((depth_extension == 1) ? 18 : 4) :
                            (width_a == 36) ? ((depth_extension == 1) ? 36: 9) :
                            (width_a == 72) ? 18 : 18;
                            
    parameter width_b_5k =  (width_b == 1) ? 1 : 
                            (width_b == 2) ? 2 :
                            (width_b == 4) ? ((depth_extension == 1) ? 4 : 1) :
                            (width_b == 9) ? ((depth_extension == 1) ? 9 : 2) :
                            (width_b == 18) ? ((depth_extension == 1) ? 18 : 4) :
                            (width_b == 36) ? ((depth_extension == 1) ? 36: 9) :
                            (width_b == 72) ? 18 : 18;

                            
    localparam [3:0] modea_sel = (width_a_5k == 1) ? 4'b1111 : 
                           (width_a_5k == 2) ? 4'b1110 :
                           (width_a_5k == 4) ? 4'b1100 :
                           (width_a_5k == 9) ? 4'b1000 :
                           (width_a_5k == 18) ? 4'b0000 : 4'b0000;
                           
    localparam [3:0] modeb_sel = (width_b_5k == 1) ? 4'b1111 : 
                           (width_b_5k == 2) ? 4'b1110 :
                           (width_b_5k == 4) ? 4'b1100 :
                           (width_b_5k == 9) ? 4'b1000 :
                           (width_b_5k == 18) ? 4'b0000 : 4'b0000;

    localparam [1:0] modea_wr = (writemode_a == "write_first") ? 2'b01 :
                          (writemode_a == "no_change") ? 2'b00 :
                          (writemode_a == "read_first") ? 2'b11 : 2'b01;
                          
    localparam [1:0] modeb_wr = (writemode_b == "write_first") ? 2'b01 :
                          (writemode_b == "no_change") ? 2'b00 :
                          (writemode_b == "read_first") ? 2'b11 : 2'b01;
                          
                            
    wire [17:0] dataina_bnk1 = (width_a_5k == 18) ? ((depth_extension == 1'b1) ? {dipa[1:0], dia[15:0]}:
                                                      (width_a_5k <= width_b_5k) ? {dipa[1:0], dia[15:0]}:
                                                      (width_b_5k == 1) ? {dipa[4],dipa[0],dia[60], dia[56], dia[52], dia[48], dia[44], dia[40], dia[36], dia[32],dia[28], dia[24], dia[20], dia[16], dia[12], dia[8], dia[4], dia[0]}:
                                                      (width_b_5k == 2) ? {dipa[4],dipa[0],dia[57:56],dia[49:48],dia[41:40],dia[33:32],dia[25:24],dia[17:16],dia[9:8],dia[1:0]}:
                                                      (width_b_5k == 4) ? {dipa[4],dipa[0],dia[51:48],dia[35:32],dia[19:16],dia[3:0]}:
                                                      (width_b_5k == 9) ? {dipa[4],dipa[0], dia[39:32], dia[7:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (width_a_5k == 9) ? ((depth_extension == 1'b1) ? {dipa[0], dipa[0], dia[7:0], dia[7:0]} :
                                                      (width_a_5k <= width_b_5k) ? {dipa[0], dipa[0], dia[7:0], dia[7:0]} :
                                                      (width_b_5k == 1) ? {dipa[0],dipa[0],dia[28], dia[24], dia[20], dia[16], dia[12], dia[8], dia[4], dia[0],dia[28], dia[24], dia[20], dia[16], dia[12], dia[8], dia[4], dia[0]}:
                                                      (width_b_5k == 2) ? {dipa[0],dipa[0],dia[25:24],dia[17:16],dia[9:8],dia[1:0],dia[25:24],dia[17:16],dia[9:8],dia[1:0]}:
                                                      (width_b_5k == 4) ? {dipa[0],dipa[0],dia[19:16],dia[3:0],dia[19:16],dia[3:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (width_a_5k == 4) ? ((depth_extension == 1'b1) ? {1'bx, 1'bx, {4{dia[3:0]}}} :
                                                      (width_a_5k <= width_b_5k) ? {1'bx, 1'bx, {4{dia[3:0]}}} :
                                                      (width_b_5k == 1) ? {1'bx, 1'bx, {4{dia[12], dia[8], dia[4], dia[0]}}}:
                                                      (width_b_5k == 2) ? {1'bx, 1'bx, {4{dia[9:8],dia[1:0]}}}:
                                                      18'bxxxxxxxxxxxxxxxxxx):
                               (width_a_5k == 2) ? {1'bx, 1'bx, {8{dia[1:0]}}} :
                               (width_a_5k == 1) ? {1'bx, 1'bx, {16{dia[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;


    wire [17:0] dataina_bnk2 = (width_a_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[3:2], dia[31:16]}:
                                                      (width_b_5k == 1) ? {dipa[5],dipa[1],dia[61], dia[57], dia[53], dia[49], dia[45], dia[41], dia[37], dia[33],dia[29], dia[25], dia[21], dia[17], dia[13], dia[9], dia[5], dia[1]}:
                                                      (width_b_5k == 2) ? {dipa[5],dipa[1],dia[59:58],dia[51:50],dia[43:42],dia[35:34],dia[27:26],dia[19:18],dia[11:10],dia[3:2]}:
                                                      (width_b_5k == 4) ? {dipa[5],dipa[1],dia[55:52],dia[39:36],dia[23:20],dia[7:4]}:
                                                      (width_b_5k == 9) ? {dipa[5],dipa[1], dia[47:40], dia[15:8]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_a_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[1], dipa[1], dia[15:8], dia[15:8]} :
                                                      (width_b_5k == 1) ? {dipa[1],dipa[1],dia[29], dia[25], dia[21], dia[17], dia[13], dia[9], dia[5], dia[1],dia[29], dia[25], dia[21], dia[17], dia[13], dia[9], dia[5], dia[1]}:
                                                      (width_b_5k == 2) ? {dipa[1],dipa[1],dia[27:26],dia[19:18],dia[11:10],dia[3:2],dia[27:26],dia[19:18],dia[11:10],dia[3:2]}:
                                                      (width_b_5k == 4) ? {dipa[1],dipa[1],dia[23:20],dia[7:4],dia[23:20],dia[7:4]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_a_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {1'bx, 1'bx, {4{dia[7:4]}}} :
                                                      (width_b_5k == 1) ? {1'bx, 1'bx, {4{ dia[13], dia[9], dia[5], dia[1]}}}:
                                                      (width_b_5k == 2) ? {1'bx, 1'bx, {4{dia[11:10],dia[3:2]}}}:18'bxxxxxxxxxxxxxxxxxx ) :
                               (width_a_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dia[3:2]}}}) :
                               (width_a_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dia[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                        
                        
   wire [17:0] dataina_bnk3 = (width_a_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[5:4], dia[47:32]}:
                                                      (width_b_5k == 1) ? {dipa[6],dipa[2],dia[62], dia[58], dia[54], dia[50], dia[46], dia[42], dia[38], dia[34],dia[30], dia[26], dia[22], dia[18], dia[14], dia[10], dia[6], dia[2]}:
                                                      (width_b_5k == 2) ? {dipa[6],dipa[2],dia[61:60],dia[53:52],dia[45:44],dia[37:36],dia[29:28],dia[21:20],dia[13:12],dia[5:4]}:
                                                      (width_b_5k == 4) ? {dipa[6],dipa[2],dia[59:56],dia[43:40],dia[27:24],dia[11:8]}:
                                                      (width_b_5k == 9) ? {dipa[6],dipa[2], dia[55:48], dia[23:16]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_a_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[2], dipa[2], dia[23:16], dia[23:16]} :
                                                      (width_b_5k == 1) ? {dipa[2],dipa[2],dia[30], dia[26], dia[22], dia[18], dia[14], dia[10], dia[6], dia[2],dia[30], dia[26], dia[22], dia[18], dia[14], dia[10], dia[6], dia[2]}:
                                                      (width_b_5k == 2) ? {dipa[2],dipa[2],dia[29:28],dia[21:20],dia[13:12],dia[5:4],dia[29:28],dia[21:20],dia[13:12],dia[5:4]}:
                                                      (width_b_5k == 4) ? {dipa[2],dipa[2],dia[27:24],dia[11:8],dia[27:24],dia[11:8]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_a_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {1'bx, 1'bx, {4{dia[11:8]}}}:
                                                      (width_b_5k == 1) ? {1'bx, 1'bx, {4{dia[14], dia[10], dia[6], dia[2]}}}:
                                                      (width_b_5k == 2) ? {1'bx, 1'bx, {4{dia[13:12],dia[5:4]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (width_a_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dia[5:4]}}}) :
                               (width_a_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dia[2]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                            
   wire [17:0] dataina_bnk4 = (width_a_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[7:6], dia[63:48]}:
                                                      (width_b_5k == 1) ? {dipa[7],dipa[3],dia[63], dia[59], dia[55], dia[51], dia[47], dia[43], dia[39], dia[35],dia[31], dia[27], dia[23], dia[19], dia[15], dia[11], dia[7], dia[3]}:
                                                      (width_b_5k == 2) ? {dipa[7],dipa[3],dia[63:62],dia[55:54],dia[47:46],dia[39:38],dia[31:30],dia[23:22],dia[15:14],dia[7:6]}:
                                                      (width_b_5k == 4) ? {dipa[7],dipa[3],dia[63:60],dia[47:44],dia[31:28],dia[15:12]}:
                                                      (width_b_5k == 9) ? {dipa[7],dipa[3], dia[63:56], dia[31:24]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_a_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {dipa[3], dipa[3], dia[31:24], dia[31:24]} :
                                                      (width_b_5k == 1) ? {dipa[3],dipa[3],dia[31], dia[27], dia[23], dia[19], dia[15], dia[11], dia[7], dia[3],dia[31], dia[27], dia[23], dia[19], dia[15], dia[11], dia[7], dia[3]}:
                                                      (width_b_5k == 2) ? {dipa[3],dipa[3],dia[31:30],dia[23:22],dia[15:14],dia[7:6],dia[31:30],dia[23:22],dia[15:14],dia[7:6]}:
                                                      (width_b_5k == 4) ? {dipa[3],dipa[3],dia[31:28],dia[15:12],dia[31:28],dia[15:12]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_a_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_a_5k <= width_b_5k) ? {1'bx, 1'bx, {4{dia[15:12]}}}:
                                                      (width_b_5k == 1) ? {1'bx, 1'bx, {4{dia[15], dia[11], dia[7], dia[3]}}}:
                                                      (width_b_5k == 2) ? {1'bx, 1'bx, {4{dia[15:14],dia[7:6]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (width_a_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dia[7:6]}}}) :
                               (width_a_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dia[3]}}}) : 18'bxxxxxxxxxxxxxxxxxx;

                
    wire [17:0] datainb_bnk1 = (width_b_5k == 18) ? ((depth_extension == 1'b1) ? {dipb[1:0], dib[15:0]}:
                                                      (width_b_5k <= width_a_5k) ? {dipb[1:0], dib[15:0]}:
                                                      (width_a_5k == 1) ? {dipb[4],dipb[0],dib[60], dib[56], dib[52], dib[48], dib[44], dib[40], dib[36], dib[32],dib[28], dib[24], dib[20], dib[16], dib[12], dib[8], dib[4], dib[0]}:
                                                      (width_a_5k == 2) ? {dipb[4],dipb[0],dib[57:56],dib[49:48],dib[41:40],dib[33:32],dib[25:24],dib[17:16],dib[9:8],dib[1:0]}:
                                                      (width_a_5k == 4) ? {dipb[4],dipb[0],dib[51:48],dib[35:32],dib[19:16],dib[3:0]}:
                                                      (width_a_5k == 9) ? {dipb[4],dipb[0], dib[39:32], dib[7:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (width_b_5k == 9) ? ((depth_extension == 1'b1) ? {dipb[0], dipb[0], dib[7:0], dib[7:0]} :
                                                      (width_b_5k <= width_a_5k) ? {dipb[0], dipb[0], dib[7:0], dib[7:0]} :
                                                      (width_a_5k == 1) ? {dipb[0],dipb[0],dib[28], dib[24], dib[20], dib[16], dib[12], dib[8], dib[4], dib[0],dib[28], dib[24], dib[20], dib[16], dib[12], dib[8], dib[4], dib[0]}:
                                                      (width_a_5k == 2) ? {dipb[0],dipb[0],dib[25:24],dib[17:16],dib[9:8],dib[1:0],dib[25:24],dib[17:16],dib[9:8],dib[1:0]}:
                                                      (width_a_5k == 4) ? {dipb[0],dipb[0],dib[19:16],dib[3:0],dib[19:16],dib[3:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (width_b_5k == 4) ? ((depth_extension == 1'b1) ? {1'bx, 1'bx, {4{dib[3:0]}}} :
                                                      (width_b_5k <= width_a_5k) ? {1'bx, 1'bx, {4{dib[3:0]}}} :
                                                      (width_a_5k == 1) ? {1'bx, 1'bx, {4{dib[12], dib[8], dib[4], dib[0]}}}:
                                                      (width_a_5k == 2) ? {1'bx, 1'bx, {4{dib[9:8],dib[1:0]}}} :18'bxxxxxxxxxxxxxxxxxx): 
                                                      
                               (width_b_5k == 2) ? {1'bx, 1'bx, {8{dib[1:0]}}} :
                               (width_b_5k == 1) ? {1'bx, 1'bx, {16{dib[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;


    wire [17:0] datainb_bnk2 = (width_b_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[3:2], dib[31:16]}:
                                                      (width_a_5k == 1) ? {dipb[5],dipb[1],dib[61], dib[57], dib[53], dib[49], dib[45], dib[41], dib[37], dib[33],dib[29], dib[25], dib[21], dib[17], dib[13], dib[9], dib[5], dib[1]}:
                                                      (width_a_5k == 2) ? {dipb[5],dipb[1],dib[59:58],dib[51:50],dib[43:42],dib[35:34],dib[27:26],dib[19:18],dib[11:10],dib[3:2]}:
                                                      (width_a_5k == 4) ? {dipb[5],dipb[1],dib[55:52],dib[39:36],dib[23:20],dib[7:4]}:
                                                      (width_a_5k == 9) ? {dipb[5],dipb[1], dib[47:40], dib[15:8]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_b_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[1], dipb[1], dib[15:8], dib[15:8]} :
                                                      (width_a_5k == 1) ? {dipb[1],dipb[1],dib[29], dib[25], dib[21], dib[17], dib[13], dib[9], dib[5], dib[1],dib[29], dib[25], dib[21], dib[17], dib[13], dib[9], dib[5], dib[1]}:
                                                      (width_a_5k == 2) ? {dipb[1],dipb[1],dib[27:26],dib[19:18],dib[11:10],dib[3:2],dib[27:26],dib[19:18],dib[11:10],dib[3:2]}:
                                                      (width_a_5k == 4) ? {dipb[1],dipb[1],dib[23:20],dib[7:4],dib[23:20],dib[7:4]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {1'bx, 1'bx, {4{dib[7:4]}}}: 
                                                      (width_a_5k == 1) ? {1'bx, 1'bx,{4{dib[13], dib[9], dib[5], dib[1]}}}:
                                                      (width_a_5k == 2) ? {1'bx, 1'bx,{4{dib[11:10],dib[3:2]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dib[3:2]}}}) :
                               (width_b_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dib[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                        
                        
   wire [17:0] datainb_bnk3 = (width_b_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[5:4], dib[47:32]}:
                                                      (width_a_5k == 1) ? {dipb[6],dipb[2],dib[62], dib[58], dib[54], dib[50], dib[46], dib[42], dib[38], dib[34],dib[30], dib[26], dib[22], dib[18], dib[14], dib[10], dib[6], dib[2]}:
                                                      (width_a_5k == 2) ? {dipb[6],dipb[2],dib[61:60],dib[53:52],dib[45:44],dib[37:36],dib[29:28],dib[21:20],dib[13:12],dib[5:4]}:
                                                      (width_a_5k == 4) ? {dipb[6],dipb[2],dib[59:56],dib[43:40],dib[27:24],dib[11:8]}:
                                                      (width_a_5k == 9) ? {dipb[6],dipb[2], dib[55:48], dib[23:16]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_b_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[2], dipb[2], dib[23:16], dib[23:16]} :
                                                      (width_a_5k == 1) ? {dipb[2],dipb[2],dib[30], dib[26], dib[22], dib[18], dib[14], dib[10], dib[6], dib[2],dib[30], dib[26], dib[22], dib[18], dib[14], dib[10], dib[6], dib[2]}:
                                                      (width_a_5k == 2) ? {dipb[2],dipb[2],dib[29:28],dib[21:20],dib[13:12],dib[5:4],dib[29:28],dib[21:20],dib[13:12],dib[5:4]}:
                                                      (width_a_5k == 4) ? {dipb[2],dipb[2],dib[27:24],dib[11:8],dib[27:24],dib[11:8]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {1'bx, 1'bx, {4{dib[11:8]}}} :
                                                      (width_a_5k == 1) ? {1'bx, 1'bx, {4{dib[14], dib[10], dib[6], dib[2]}}}:
                                                      (width_a_5k == 2) ? {1'bx, 1'bx, {4{dib[13:12],dib[5:4]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dib[5:4]}}}) :
                               (width_b_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dib[2]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                            
   wire [17:0] datainb_bnk4 = (width_b_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[7:6], dib[63:48]}:
                                                      (width_a_5k == 1) ? {dipb[7],dipb[3],dib[63], dib[59], dib[55], dib[51], dib[47], dib[43], dib[39], dib[35],dib[31], dib[27], dib[23], dib[19], dib[15], dib[11], dib[7], dib[3]}:
                                                      (width_a_5k == 2) ? {dipb[7],dipb[3],dib[63:62],dib[55:54],dib[47:46],dib[39:38],dib[31:30],dib[23:22],dib[15:14],dib[7:6]}:
                                                      (width_a_5k == 4) ? {dipb[7],dipb[3],dib[63:60],dib[47:44],dib[31:28],dib[15:12]}:
                                                      (width_a_5k == 9) ? {dipb[7],dipb[3], dib[63:56], dib[31:24]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (width_b_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {dipb[3], dipb[3], dib[31:24], dib[31:24]} :
                                                      (width_a_5k == 1) ? {dipb[3],dipb[3],dib[31], dib[27], dib[23], dib[19], dib[15], dib[11], dib[7], dib[3],dib[31], dib[27], dib[23], dib[19], dib[15], dib[11], dib[7], dib[3]}:
                                                      (width_a_5k == 2) ? {dipb[3],dipb[3],dib[31:30],dib[23:22],dib[15:14],dib[7:6],dib[31:30],dib[23:22],dib[15:14],dib[7:6]}:
                                                      (width_a_5k == 4) ? {dipb[3],dipb[3],dib[31:28],dib[15:12],dib[31:28],dib[15:12]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (width_b_5k <= width_a_5k) ? {1'bx, 1'bx, {4{dib[15:12]}}} :
                                                      (width_a_5k == 1) ? {1'bx, 1'bx, {4{dib[15], dib[11], dib[7], dib[3]}}}:
                                                      (width_a_5k == 2) ? {1'bx, 1'bx, {4{dib[15:14],dib[7:6]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (width_b_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{dib[7:6]}}}) :
                               (width_b_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{dib[3]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                            
                            
    wire [7:0] dopa_buf0;
    wire [3:0] dopb_buf0;
    
    wire [7:0] dopa_buf1;
    wire [3:0] dopb_buf1;
    
    integer i;
    
    // assign dopa =   (depth_extension == 1'b1) ? dopa_buf1 :
                    // (width_a_5k <= width_b_5k) ? dopa_buf1 :
                    // (width_b_5k == 9) ? {dopa_buf1[7], dopa_buf1[5], dopa_buf1[3], dopa_buf1[1], 
                                        // dopa_buf1[6], dopa_buf1[4], dopa_buf1[2], dopa_buf1[0]} : dopa_buf1;
    assign dopa = dopa_buf1;                      
    assign dopb = dopb_buf1; 
    
    assign dopa_buf1 =  (depth_extension == 1'b1) ? dopa_buf0 :
                        (width_a_5k <= width_b_5k) ? dopa_buf0 :
                        (width_b_5k == 9) ? {dopa_buf0[7], dopa_buf0[5], dopa_buf0[3], dopa_buf0[1], 
                                            dopa_buf0[6], dopa_buf0[4], dopa_buf0[2], dopa_buf0[0]} : dopa_buf0;
                          
    assign dopb_buf1 =  dopb_buf0;    
                                                                                    
    wire [17:0] dataout_bnk1;
    wire [17:0] dataout_bnk2;
    wire [17:0] dataout_bnk3;
    wire [17:0] dataout_bnk4;

    assign dopb_buf0 =  (depth_extension == 1'b1) ? {3'bxxx, dataout_bnk1[17]} : 
                        (depth_extension == 1'b1) ? {2'bxx, dataout_bnk3[17], dataout_bnk1[17]} : 
                        {dataout_bnk4[17], dataout_bnk3[17], dataout_bnk2[17], dataout_bnk1[17]};
                 
    assign dopa_buf0[7:4] = (depth_extension == 1'b1) ? 4'bxxxx : 
                            (depth_extension == 1'b1) ? 4'bxxxx : 
                            (width_a_5k == 18) ?    {dataout_bnk4[17], dataout_bnk4[16], dataout_bnk3[17], dataout_bnk3[16]}
                                                    :4'bxxxx;

    assign dopa_buf0[3:2] = (depth_extension == 1'b1) ? 2'bxx : 
                            (depth_extension == 1'b1) ? ((width_a_5k == 18) ? {dataout_bnk3[17], dataout_bnk3[16]} : 
                                                                                2'bxx) : 
                            (width_a_5k == 18) ?    {dataout_bnk2[17], dataout_bnk2[16]} : 
                                                    {dataout_bnk4[8], dataout_bnk3[8]};

    assign dopa_buf0[1:0] = (depth_extension == 1'b1) ? ((width_a_5k == 18) ? {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                                                {1'bx, dataout_bnk1[8]}) : 
                            (depth_extension == 1'b1) ? ((width_a_5k == 18) ? {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                                                {dataout_bnk3[8], dataout_bnk1[8]}) : 
                            (width_a_5k == 18) ?    {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                    {dataout_bnk2[8], dataout_bnk1[8]};
                                                
    assign doa = width_a_5k==1 ? {60'h0,dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]} :
                 width_a_5k==2 ? {56'h0,dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]} :
                 width_a_5k==4 ? ((depth_extension == 1'b1) ? {48'h0,dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]} :
                                   (width_b_5k >= width_a_5k) ? {48'h0,dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]} :                           
                                   (width_b_5k == 2) ? {48'h0,dataout_bnk4[3:2],dataout_bnk3[3:2],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (width_b_5k == 1) ? {48'h0,dataout_bnk4[3],dataout_bnk3[3],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk4[2],dataout_bnk3[2],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk4[1],dataout_bnk3[1],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]}: 
                                   {48'h0,dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]}):
                                   
                 width_a_5k==9 ? ((depth_extension == 1'b1) ? {32'h0,dataout_bnk4[7:0],dataout_bnk3[7:0],dataout_bnk2[7:0],dataout_bnk1[7:0]} :
                                   (width_b_5k >= width_a_5k) ?{32'h0,dataout_bnk4[7:0],dataout_bnk3[7:0],dataout_bnk2[7:0],dataout_bnk1[7:0]} :                            
                                   (width_b_5k == 4) ? {dataout_bnk4[7:4],dataout_bnk3[7:4],dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (width_b_5k == 2) ? {dataout_bnk4[7:6],dataout_bnk3[7:6],dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk4[5:4],dataout_bnk3[5:4],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk4[3:2],dataout_bnk3[3:2],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (width_b_5k == 1) ? {dataout_bnk4[7],dataout_bnk3[7],dataout_bnk2[7],dataout_bnk1[7],dataout_bnk4[6],dataout_bnk3[6],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk4[5],dataout_bnk3[5],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk4[4],dataout_bnk3[4],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk4[3],dataout_bnk3[3],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk4[2],dataout_bnk3[2],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk4[1],dataout_bnk3[1],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]}:
                                   {dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0]  }) :
                 
                 width_a_5k==18 ? ((depth_extension == 1'b1) ? {dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (width_b_5k >= width_a_5k) ?{dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (width_b_5k == 9) ? {dataout_bnk4[15:8],dataout_bnk3[15:8],dataout_bnk2[15:8],dataout_bnk1[15:8],dataout_bnk4[7:0],dataout_bnk3[7:0],dataout_bnk2[7:0],dataout_bnk1[7:0]  }:
                                   (width_b_5k == 4) ? {dataout_bnk4[15:12],dataout_bnk3[15:12],dataout_bnk2[15:12],dataout_bnk1[15:12],dataout_bnk4[11:8],dataout_bnk3[11:8],dataout_bnk2[11:8],dataout_bnk1[11:8],dataout_bnk4[7:4],dataout_bnk3[7:4],dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (width_b_5k == 2) ? {dataout_bnk4[15:14],dataout_bnk3[15:14],dataout_bnk2[15:14],dataout_bnk1[15:14],dataout_bnk4[13:12],dataout_bnk3[13:12],dataout_bnk2[13:12],dataout_bnk1[13:12],dataout_bnk4[11:10],dataout_bnk3[11:10],dataout_bnk2[11:10],dataout_bnk1[11:10],dataout_bnk4[9:8],dataout_bnk3[9:8],dataout_bnk2[9:8],dataout_bnk1[9:8],dataout_bnk4[7:6],dataout_bnk3[7:6],dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk4[5:4],dataout_bnk3[5:4],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk4[3:2],dataout_bnk3[3:2],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (width_b_5k == 1) ? {dataout_bnk4[15],dataout_bnk3[15],dataout_bnk2[15],dataout_bnk1[15],dataout_bnk4[14],dataout_bnk3[14],dataout_bnk2[14],dataout_bnk1[14],dataout_bnk4[13],dataout_bnk3[13],dataout_bnk2[13],dataout_bnk1[13],dataout_bnk4[12],dataout_bnk3[12],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk4[11],dataout_bnk3[11],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk4[10],dataout_bnk3[10],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk4[9],dataout_bnk3[9],dataout_bnk2[9],dataout_bnk1[9],dataout_bnk4[8],dataout_bnk3[8],dataout_bnk2[8],dataout_bnk1[8],dataout_bnk4[7],dataout_bnk3[7],dataout_bnk2[7],dataout_bnk1[7],dataout_bnk4[6],dataout_bnk3[6],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk4[5],dataout_bnk3[5],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk4[4],dataout_bnk3[4],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk4[3],dataout_bnk3[3],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk4[2],dataout_bnk3[2],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk4[1],dataout_bnk3[1],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]}:{dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0] }) :
                 64'hxxxx_xxxx_xxxx_xxxx;             
                 
    assign dob = width_b_5k==1 ? {28'h0,dataout_bnk4[9],dataout_bnk3[9],dataout_bnk2[9],dataout_bnk1[9]} :
                 width_b_5k==2 ? {24'h0,dataout_bnk4[10:9],dataout_bnk3[10:9],dataout_bnk2[10:9],dataout_bnk1[10:9]} :
                 width_b_5k==4 ? ((depth_extension == 1'b1) ? {16'h0,dataout_bnk4[12:9],dataout_bnk3[12:9],dataout_bnk2[12:9],dataout_bnk1[12:9]} :
                                   (width_a_5k >= width_b_5k) ? {16'h0,dataout_bnk4[12:9],dataout_bnk3[12:9],dataout_bnk2[12:9],dataout_bnk1[12:9]} :                            
                                   (width_a_5k == 2) ? {16'h0,dataout_bnk4[12:11],dataout_bnk3[12:11],dataout_bnk2[12:11],dataout_bnk1[12:11],dataout_bnk4[10:9],dataout_bnk3[10:9],dataout_bnk2[10:9],dataout_bnk1[10:9]}:
                                   (width_a_5k == 1) ? {16'h0,dataout_bnk4[12],dataout_bnk3[12],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk4[11],dataout_bnk3[11],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk4[10],dataout_bnk3[10],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk4[9],dataout_bnk3[9],dataout_bnk2[9],dataout_bnk1[9]}:
                                   {16'h0,dataout_bnk4[12:9],dataout_bnk3[12:9],dataout_bnk2[12:9],dataout_bnk1[12:9]}) :
                                   
                 width_b_5k==9 ? ((depth_extension == 1'b1) ? {dataout_bnk4[16:9],dataout_bnk3[16:9],dataout_bnk2[16:9],dataout_bnk1[16:9]} :
                                   (width_a_5k >= width_b_5k) ?{dataout_bnk4[16:9],dataout_bnk3[16:9],dataout_bnk2[16:9],dataout_bnk1[16:9]} :                            
                                   (width_a_5k == 4) ? {dataout_bnk4[16:13],dataout_bnk3[16:13],dataout_bnk2[16:13],dataout_bnk1[16:13],dataout_bnk4[12:9],dataout_bnk3[12:9],dataout_bnk2[12:9],dataout_bnk1[12:9]  }:
                                   (width_a_5k == 2) ? {dataout_bnk4[16:15],dataout_bnk3[16:15],dataout_bnk2[16:15],dataout_bnk1[16:15],dataout_bnk4[14:13],dataout_bnk3[14:13],dataout_bnk2[14:13],dataout_bnk1[14:13],dataout_bnk4[12:11],dataout_bnk3[12:11],dataout_bnk2[12:11],dataout_bnk1[12:11],dataout_bnk4[10:9],dataout_bnk3[10:9],dataout_bnk2[10:9],dataout_bnk1[10:9]}:
                                   (width_a_5k == 1) ? {dataout_bnk4[16],dataout_bnk3[16],dataout_bnk2[16],dataout_bnk1[16],dataout_bnk4[15],dataout_bnk3[15],dataout_bnk2[15],dataout_bnk1[15],dataout_bnk4[14],dataout_bnk3[14],dataout_bnk2[14],dataout_bnk1[14],dataout_bnk4[13],dataout_bnk3[13],dataout_bnk2[13],dataout_bnk1[13],dataout_bnk4[12],dataout_bnk3[12],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk4[11],dataout_bnk3[11],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk4[10],dataout_bnk3[10],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk4[9],dataout_bnk3[9],dataout_bnk2[9],dataout_bnk1[9]}:
                                   {dataout_bnk4[16:9],dataout_bnk3[16:9],dataout_bnk2[16:9],dataout_bnk1[16:9]}) :
                 32'hxxxx_xxxx;
    wire [1:0] regen = (rammode == "tdp") ? {regceb, regcea} : {regcea, regcea};
    
    // address translation
               
    //sp mode
    localparam sp_addr_lbit =  (width_a == 1) ? 0 : (width_a == 2) ? 1 : 
                               (width_a == 4) ? 2 : (width_a == 9) ? 3 : 
                               (width_a == 18) ? 4 : (width_a == 36) ? 3 : 
                               (width_a == 72) ? 4: 0; 
 
    //sdp mode 
    localparam sdp_raddr_lbit = (width_a == 1) ? 0 :
                                (width_a == 2) ? 1 : 
                                (width_a == 4) ? ((width_b == 36 || width_b == 72) ? 0 : 2) : 
                                (width_a == 9) ? ((width_b == 36 || width_b == 72) ? 1 : 3) : 
                                (width_a == 18) ? ((width_b == 36 || width_b == 72) ? 2 : 4) : 
                                (width_a == 36) ? 3 :
                                (width_a == 72) ? 4 : 0;
                       
    localparam sdp_waddr_lbit = (width_b == 1) ? 0 :
                                (width_b == 2) ? 1 : 
                                (width_b == 4) ? ((width_a == 36 || width_a == 72) ? 0 : 2) : 
                                (width_b == 9) ? ((width_a == 36 || width_a == 72) ? 1 : 3) : 
                                (width_b == 18) ? ((width_a == 36 || width_a == 72) ? 2 : 4) : 
                                (width_b == 36) ? 3 : 
                                (width_b == 72) ? 4: 0;
    //tdp mode
    localparam tdp_addra_lbit = (width_a == 1) ? 0 : 
                                (width_a == 2) ? 1 : 
                                (width_a == 4) ? ((width_b== 18 ||width_b == 36) ? 0:2) : 
                                (width_a == 9) ? ((width_b== 18 ||width_b == 36) ? 1:3) : 
                                (width_a == 18) ? 2 :
                                (width_a == 36) ? 3 : 0;
                   
    localparam tdp_addrb_lbit = (width_b == 1) ? 0 : (width_b == 2) ? 1 : 
                                (width_b == 4) ? ((width_a== 18 ||width_a == 36) ? 0:2) : 
                                (width_b == 9) ? ((width_a== 18 ||width_a == 36) ? 1:3) : 
                                (width_b == 18) ? 2 :
                                (width_b == 36) ? 3 : 0;
           
    localparam addra_lbit = (rammode == "sp")  ? sp_addr_lbit :
                            (rammode == "sdp") ? sdp_raddr_lbit :
                            (rammode == "tdp") ? tdp_addra_lbit : 0;
    localparam addrb_lbit = (rammode == "sp")  ? sp_addr_lbit :
                            (rammode == "sdp") ? sdp_waddr_lbit :
                            (rammode == "tdp") ? tdp_addrb_lbit : 0;
    //translation
    wire [13:0] addra_input;
    wire [13:0] addrb_input;
    
    localparam  addr_width_a = (width_a == 1)  ? 14 : (width_a == 2)  ? 13 :
                               (width_a == 4)  ? 12 : (width_a == 8)  ? 11 :
                               (width_a == 9)  ? 11 : (width_a == 16) ? 10 :
                               (width_a == 18) ? 10 : (width_a == 32) ? 9 :
                               (width_a == 36) ? 9  : (width_a == 64) ? 8 :
                               (width_a == 72) ? 8  :0;
    localparam  addr_width_b = (width_b == 1)  ? 14 : (width_b == 2)  ? 13 :
                               (width_b == 4)  ? 12 : (width_b == 8)  ? 11 :
                               (width_b == 9)  ? 11 : (width_b == 16) ? 10 :
                               (width_b == 18) ? 10 : (width_b == 32) ? 9 :
                               (width_b == 36) ? 9  : (width_b == 64) ? 8 :
                               (width_b == 72) ? 8  : 1;//sp mode not use port b default 1 for addrb_input[addrb_lbit + addr_width_b - 1 : addrb_lbit] = addrb; when with_b=0
                               
    assign addra_input[addra_lbit + addr_width_a - 1 : addra_lbit] = addra;    
    if (addra_lbit > 0)
        assign addra_input[addra_lbit - 1 : 0] = 0;
    if (addra_lbit + addr_width_a < 14)
        assign addra_input[13 : addra_lbit + addr_width_a] = 0;
        
    assign addrb_input[addrb_lbit + addr_width_b - 1 : addrb_lbit] = addrb;
    if (addrb_lbit > 0)
        assign addrb_input[addrb_lbit - 1 : 0] = 0;
    if (addrb_lbit + addr_width_b < 14)
        assign addrb_input[13 : addrb_lbit + addr_width_b] = 0; 
    
BRAM18KV1 # (
    .DEPTH_EXT_MODE23        (depth_extension),
    .DEPTH_EXT_MODE01        (depth_extension),
    .ECC_DEC_EN                (eccreaden),
    .ECC_ENC_EN                (eccwriteen),
    
    .EMB5K_4_MODEA_SEL      (modea_sel),
    .EMB5K_4_MODEB_SEL      (modeb_sel),
    .EMB5K_4_PORTA_BYPASS   (1'b0),
    .EMB5K_4_PORTA_CE       (1'b1),
    .EMB5K_4_PORTA_REG_OUT  (outreg_a),
    .EMB5K_4_PORTA_WR_MODE  (modea_wr),
    .EMB5K_4_PORTA_CKINV    (clka_inv),
    .EMB5K_4_PORTB_BYPASS   (1'b0),
    .EMB5K_4_PORTB_CE       (1'b1),
    .EMB5K_4_PORTB_REG_OUT  (outreg_b),
    .EMB5K_4_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_4_PORTB_CKINV    (clkb_inv),
    
    .EMB5K_3_MODEA_SEL      (modea_sel),
    .EMB5K_3_MODEB_SEL      (modeb_sel),
    .EMB5K_3_PORTA_BYPASS   (1'b0),
    .EMB5K_3_PORTA_CE       (1'b1),
    .EMB5K_3_PORTA_REG_OUT  (outreg_a),
    .EMB5K_3_PORTA_WR_MODE  (modea_wr),
    .EMB5K_3_PORTA_CKINV    (clka_inv),
    .EMB5K_3_PORTB_BYPASS   (1'b0),
    .EMB5K_3_PORTB_CE       (1'b1),
    .EMB5K_3_PORTB_REG_OUT  (outreg_b),
    .EMB5K_3_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_3_PORTB_CKINV    (clkb_inv),
    
    .EMB5K_2_MODEA_SEL      (modea_sel),
    .EMB5K_2_MODEB_SEL      (modeb_sel),
    .EMB5K_2_PORTA_BYPASS   (1'b0),
    .EMB5K_2_PORTA_CE       (1'b1),
    .EMB5K_2_PORTA_REG_OUT  (outreg_a),
    .EMB5K_2_PORTA_WR_MODE  (modea_wr),
    .EMB5K_2_PORTA_CKINV    (clka_inv),
    .EMB5K_2_PORTB_BYPASS   (1'b0),
    .EMB5K_2_PORTB_CE       (1'b1),
    .EMB5K_2_PORTB_REG_OUT  (outreg_b),
    .EMB5K_2_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_2_PORTB_CKINV    (clkb_inv),
    
    .EMB5K_1_MODEA_SEL      (modea_sel),
    .EMB5K_1_MODEB_SEL      (modeb_sel),
    .EMB5K_1_PORTA_BYPASS   (1'b0),
    .EMB5K_1_PORTA_CE       (1'b1),
    .EMB5K_1_PORTA_REG_OUT  (outreg_a),
    .EMB5K_1_PORTA_WR_MODE  (modea_wr),
    .EMB5K_1_PORTA_CKINV    (clka_inv),
    .EMB5K_1_PORTB_BYPASS   (1'b0),
    .EMB5K_1_PORTB_CE       (1'b1),
    .EMB5K_1_PORTB_REG_OUT  (outreg_b),
    .EMB5K_1_PORTB_WR_MODE  (modeb_wr),
    .EMB5K_1_PORTB_CKINV    (clkb_inv),
    
    .EXT_18K                (extension18k),
    .FIFO_EN                (1'b0),
    .PORTA_PROG             (8'b11110000),
    .PORTB_PROG             (8'b00001111),
    .WIDTH_EXT_MODE23       (width_extension),
    .WIDTH_EXT_MODE01       (width_extension)
)

u0_emb18k_core (
    .a_addr_ext                ({addra_input[13], addra_input[12]}),
    .b_addr_ext                ({addrb_input[13], addrb_input[12]}),
    
    .c1r4_aa                (addra_input[11:0]),
    .c1r4_ab                (addrb_input[11:0]),
    .c1r4_cea                (cea),
    .c1r4_ceb                (ceb),
    .c1r4_clka                (clka),
    .c1r4_clkb                (clkb),
    .c1r4_da                (dataina_bnk4),
    .c1r4_db                (datainb_bnk4),
    .c1r4_rstna                (regsra),
    .c1r4_rstnb                (regsrb),
    .c1r4_wea                (wea[3]),
    .c1r4_web                (web[3]),
    .c1r4_user_ena          (regen[0]),
    .c1r4_user_enb          (regen[1]), 
     
    .c1r3_aa                (addra_input[11:0]),
    .c1r3_ab                (addrb_input[11:0]),
    .c1r3_cea                (cea),
    .c1r3_ceb                (ceb),
    .c1r3_clka                (clka),
    .c1r3_clkb                (clkb),
    .c1r3_da                (dataina_bnk3),
    .c1r3_db                (datainb_bnk3),
    .c1r3_rstna                (regsra),
    .c1r3_rstnb                (regsrb),
    .c1r3_wea                (wea[2]),
    .c1r3_web                (web[2]),
    .c1r3_user_ena          (regen[0]),
    .c1r3_user_enb          (regen[1]), 
     
    .c1r2_aa                (addra_input[11:0]),
    .c1r2_ab                (addrb_input[11:0]),
    .c1r2_cea                (cea),
    .c1r2_ceb                (ceb),
    .c1r2_clka                (clka),
    .c1r2_clkb                (clkb),
    .c1r2_da                (dataina_bnk2),
    .c1r2_db                (datainb_bnk2),
    .c1r2_rstna                (regsra),
    .c1r2_rstnb                (regsrb),
    .c1r2_wea                (wea[1]),
    .c1r2_web                (web[1]),
    .c1r2_user_ena          (regen[0]),
    .c1r2_user_enb          (regen[1]), 
    
    .c1r1_aa                (addra_input[11:0]),
    .c1r1_ab                (addrb_input[11:0]),
    .c1r1_cea                (cea),
    .c1r1_ceb                (ceb),
    .c1r1_clka                (clka),
    .c1r1_clkb                (clkb),
    .c1r1_da                (dataina_bnk1),
    .c1r1_db                (datainb_bnk1),
    .c1r1_rstna                (regsra),
    .c1r1_rstnb                (regsrb),
    .c1r1_wea                (wea[0]),
    .c1r1_web                (web[0]),
    .c1r1_user_ena          (regen[0]),
    .c1r1_user_enb          (regen[1]),   
 
    .rd_mem_n                (1'b0),
    .rptr                    (14'b0),
    .wptr                    (14'b0),
    .wr_mem_n                (1'b0),
        
    .c1r4_q                    (dataout_bnk4),
    .c1r3_q                    (dataout_bnk3),
    .c1r2_q                    (dataout_bnk2),
    .c1r1_q                    (dataout_bnk1),
    .eccindberr             (eccindberr),
    .eccinsberr             (eccinsberr),
    .eccoutdberr            (eccoutdberr),
    .eccoutsberr            (eccoutsberr),
    .err_addr                  (eccreadaddr) 
    );



wire GSR;
glbsr inst( .GSR( GSR )) ;

initial
begin
    @(posedge GSR);
    for (i = 0; i < 16; i = i + 1)
    begin
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i    ] <= {initp_00[i*2+1   -:2 ], init_00[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+16 ] <= {initp_00[i*2+33  -:2 ], init_01[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+32 ] <= {initp_00[i*2+65  -:2 ], init_02[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+48 ] <= {initp_00[i*2+97  -:2 ], init_03[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+64 ] <= {initp_00[i*2+129 -:2 ], init_04[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+80 ] <= {initp_00[i*2+161 -:2 ], init_05[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+96 ] <= {initp_00[i*2+193 -:2 ], init_06[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+112] <= {initp_00[i*2+225 -:2 ], init_07[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+128] <= {initp_01[i*2+1   -:2 ], init_08[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+144] <= {initp_01[i*2+33  -:2 ], init_09[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+160] <= {initp_01[i*2+65  -:2 ], init_0a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+176] <= {initp_01[i*2+97  -:2 ], init_0b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+192] <= {initp_01[i*2+129 -:2 ], init_0c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+208] <= {initp_01[i*2+161 -:2 ], init_0d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+224] <= {initp_01[i*2+193 -:2 ], init_0e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_1.emb5k_top.mem[i+240] <= {initp_01[i*2+225 -:2 ], init_0f[i*16+15 -:16 ]};

        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i    ] <= {initp_02[i*2+1   -:2 ], init_10[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+16 ] <= {initp_02[i*2+33  -:2 ], init_11[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+32 ] <= {initp_02[i*2+65  -:2 ], init_12[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+48 ] <= {initp_02[i*2+97  -:2 ], init_13[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+64 ] <= {initp_02[i*2+129 -:2 ], init_14[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+80 ] <= {initp_02[i*2+161 -:2 ], init_15[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+96 ] <= {initp_02[i*2+193 -:2 ], init_16[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+112] <= {initp_02[i*2+225 -:2 ], init_17[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+128] <= {initp_03[i*2+1   -:2 ], init_18[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+144] <= {initp_03[i*2+33  -:2 ], init_19[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+160] <= {initp_03[i*2+65  -:2 ], init_1a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+176] <= {initp_03[i*2+97  -:2 ], init_1b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+192] <= {initp_03[i*2+129 -:2 ], init_1c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+208] <= {initp_03[i*2+161 -:2 ], init_1d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+224] <= {initp_03[i*2+193 -:2 ], init_1e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_2.emb5k_top.mem[i+240] <= {initp_03[i*2+225 -:2 ], init_1f[i*16+15 -:16 ]};

        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i    ] <= {initp_04[i*2+1   -:2 ], init_20[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+16 ] <= {initp_04[i*2+33  -:2 ], init_21[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+32 ] <= {initp_04[i*2+65  -:2 ], init_22[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+48 ] <= {initp_04[i*2+97  -:2 ], init_23[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+64 ] <= {initp_04[i*2+129 -:2 ], init_24[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+80 ] <= {initp_04[i*2+161 -:2 ], init_25[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+96 ] <= {initp_04[i*2+193 -:2 ], init_26[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+112] <= {initp_04[i*2+225 -:2 ], init_27[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+128] <= {initp_05[i*2+1   -:2 ], init_28[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+144] <= {initp_05[i*2+33  -:2 ], init_29[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+160] <= {initp_05[i*2+65  -:2 ], init_2a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+176] <= {initp_05[i*2+97  -:2 ], init_2b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+192] <= {initp_05[i*2+129 -:2 ], init_2c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+208] <= {initp_05[i*2+161 -:2 ], init_2d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+224] <= {initp_05[i*2+193 -:2 ], init_2e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_3.emb5k_top.mem[i+240] <= {initp_05[i*2+225 -:2 ], init_2f[i*16+15 -:16 ]};

        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i    ] <= {initp_06[i*2+1   -:2 ], init_30[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+16 ] <= {initp_06[i*2+33  -:2 ], init_31[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+32 ] <= {initp_06[i*2+65  -:2 ], init_32[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+48 ] <= {initp_06[i*2+97  -:2 ], init_33[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+64 ] <= {initp_06[i*2+129 -:2 ], init_34[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+80 ] <= {initp_06[i*2+161 -:2 ], init_35[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+96 ] <= {initp_06[i*2+193 -:2 ], init_36[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+112] <= {initp_06[i*2+225 -:2 ], init_37[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+128] <= {initp_07[i*2+1   -:2 ], init_38[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+144] <= {initp_07[i*2+33  -:2 ], init_39[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+160] <= {initp_07[i*2+65  -:2 ], init_3a[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+176] <= {initp_07[i*2+97  -:2 ], init_3b[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+192] <= {initp_07[i*2+129 -:2 ], init_3c[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+208] <= {initp_07[i*2+161 -:2 ], init_3d[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+224] <= {initp_07[i*2+193 -:2 ], init_3e[i*16+15 -:16 ]};
        u0_emb18k_core.emb5k_core_4.emb5k_top.mem[i+240] <= {initp_07[i*2+225 -:2 ], init_3f[i*16+15 -:16 ]};
    end
end
    
endmodule // EMB18K

// end of EMB18K

module FIFO5K (dout, doutp, din, dinp, writeclk, readclk, writeen, readen, reset, regce, 
            writesave, writedrop, full, empty, almostfull, almostempty, overflow, underflow, writedropflag);

    output [15:0] dout;
    output [1:0] doutp;
    output full, empty;
    output almostfull, almostempty;
    output overflow, underflow;
    output writedropflag;
    
    input [15:0] din;
    input [1:0] dinp;
    input writeclk, readclk;
    input writeen, readen;
    input reset, regce;
    input writesave, writedrop;

    parameter almostemptyth = 12'b0;
    parameter almostfullth = 12'b0;
    parameter writewidth = 1;
    parameter readwidth = 1;
    parameter outreg = 0;
    parameter peek = 1'b0;
    parameter readclk_inv = 1'b0;
    parameter writeclk_inv = 1'b0;


    parameter read_sel =    (readwidth == 1) ? 4'b1111 : 
                            (readwidth == 2) ? 4'b1110 :
                            (readwidth == 4) ? 4'b1100 :
                            (readwidth == 9) ? 4'b1000 :
                            (readwidth == 18) ? 4'b0000 : 4'bxxxx;    

    parameter write_sel =   (writewidth == 1) ? 4'b1111 : 
                            (writewidth == 2) ? 4'b1110 :
                            (writewidth == 4) ? 4'b1100 :
                            (writewidth == 9) ? 4'b1000 :
                            (writewidth == 18) ? 4'b0000 : 4'bxxxx;
                            
    parameter read_data_width = (readwidth == 1) ? 1 : 
                                (readwidth == 2) ? 2 :
                                (readwidth == 4) ? 4 :
                                (readwidth == 9) ? 8 :
                                (readwidth == 18) ? 16 : 0;
                                
    parameter write_data_width =    (writewidth == 1) ? 1 : 
                                    (writewidth == 2) ? 2 :
                                    (writewidth == 4) ? 4 :
                                    (writewidth == 9) ? 8 :
                                    (writewidth == 18) ? 16 : 0;   
                            
    parameter EXT_18K = 1'b0;
    parameter DEPTH_EXT_MODE01 = 1'b0;
    
    reg finish_error = 0;
    initial begin
        if (peek == 1'b1 && outreg == 0)
        begin
            $display("DRC Error : outreg = 0 is invalid when peek is set to 1 on FIFO5K instance %m.");
            finish_error = 1;
        end
    end
                           
    wire rd_mem_n;
    wire [13:0]	rptr;
    wire [13:0]	wptr;
    wire wr_mem_n;

    wire peek_en;
    wire peek_rd_en;
    
    wire [17:0] datain =    (writewidth == 18) ? {dinp, din} : 
                            (writewidth == 9) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                            (writewidth == 4) ? {1'bx, 1'bx, {4{din[3:0]}}} :
                            (writewidth == 2) ? {1'bx, 1'bx, {8{din[1:0]}}} :
                            (writewidth == 1) ? {1'bx, 1'bx, {16{din[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;
    
    wire [17:0] dataout;
    assign doutp[1] = dataout[17];
    assign doutp[0] = (readwidth == 18) ? dataout[16] : dataout[8];
    assign dout = dataout[15:0];
    
    parameter prog_full = (almostfullth + peek * 2) * write_data_width;
    parameter prog_empty = (almostemptyth - peek * 2) * read_data_width;
    
    reg [11:0] progemptyaddr_reg = prog_empty;
    reg [11:0] progfulladdr_reg = prog_full; 
                           
FIFOCTRL18KV1 # (
	.USR_PF		({2'b00, prog_full}),
	.USR_PE		({2'b00, prog_empty}),
	.PEEK_MODE	(peek),
	.FIFO_EN	(1'b1),
	.R_WIDTH	(read_sel),
	.W_WIDTH	(write_sel),
	.DEPTH_EXT_MODE	({EXT_18K, DEPTH_EXT_MODE01})
)

 u0_fifo_ctrl (
	.rst_n		(reset),
	.rd_req_n	(readen),
	.wr_req_n	(writeen),
	.clka		(readclk),
	.clkb		(writeclk),
	.write_drop	(writedrop),
	.write_save	(writesave),

	.full		(full),
	.empty		(empty),
	.prog_full	(almostfull),
	.prog_empty	(almostempty),
	.wptr		(wptr[13:0]),
	.rptr		(rptr[13:0]),
	.wr_mem_n	(wr_mem_n),
	.rd_mem_n	(rd_mem_n),
	.overflow	(overflow),
	.underflow	(underflow),
    .wrdp_rd_flag(writedropflag),
	.peek_en	(peek_en),
    .peek_rd_en (peek_rd_en)
);

BRAM18KV1 # (
    .DEPTH_EXT_MODE23       (1'b0),
    .DEPTH_EXT_MODE01       (1'b0),
    .ECC_DEC_EN             (1'b0),
    .ECC_ENC_EN             (1'b0),

    .EMB5K_4_MODEA_SEL      (),
    .EMB5K_4_MODEB_SEL      (),
    .EMB5K_4_PORTA_BYPASS   (),
    .EMB5K_4_PORTA_CE       (),
    .EMB5K_4_PORTA_REG_OUT  (),
    .EMB5K_4_PORTA_WR_MODE  (),
    .EMB5K_4_PORTA_CKINV    (),
    .EMB5K_4_PORTB_BYPASS   (),
    .EMB5K_4_PORTB_CE       (),
    .EMB5K_4_PORTB_REG_OUT  (),
    .EMB5K_4_PORTB_WR_MODE  (),
    .EMB5K_4_PORTB_CKINV    (),
    
    .EMB5K_3_MODEA_SEL      (),
    .EMB5K_3_MODEB_SEL      (),
    .EMB5K_3_PORTA_BYPASS   (),
    .EMB5K_3_PORTA_CE       (),
    .EMB5K_3_PORTA_REG_OUT  (),
    .EMB5K_3_PORTA_WR_MODE  (),
    .EMB5K_3_PORTA_CKINV    (),
    .EMB5K_3_PORTB_BYPASS   (),
    .EMB5K_3_PORTB_CE       (),
    .EMB5K_3_PORTB_REG_OUT  (),
    .EMB5K_3_PORTB_WR_MODE  (),
    .EMB5K_3_PORTB_CKINV    (),
    
    .EMB5K_2_MODEA_SEL      (),
    .EMB5K_2_MODEB_SEL      (),
    .EMB5K_2_PORTA_BYPASS   (),
    .EMB5K_2_PORTA_CE       (),
    .EMB5K_2_PORTA_REG_OUT  (),
    .EMB5K_2_PORTA_WR_MODE  (),
    .EMB5K_2_PORTA_CKINV    (),
    .EMB5K_2_PORTB_BYPASS   (),
    .EMB5K_2_PORTB_CE       (),
    .EMB5K_2_PORTB_REG_OUT  (),
    .EMB5K_2_PORTB_WR_MODE  (),
    .EMB5K_2_PORTB_CKINV    (),
    
    .EMB5K_1_MODEA_SEL      (read_sel),
    .EMB5K_1_MODEB_SEL      (write_sel),
    .EMB5K_1_PORTA_BYPASS   (1'b0),
    .EMB5K_1_PORTA_CE       (1'b1),
    .EMB5K_1_PORTA_REG_OUT  (outreg),
    .EMB5K_1_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_1_PORTA_CKINV    (readclk_inv),
    .EMB5K_1_PORTB_BYPASS   (1'b0),
    .EMB5K_1_PORTB_CE       (1'b1),
    .EMB5K_1_PORTB_REG_OUT  (outreg),
    .EMB5K_1_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_1_PORTB_CKINV    (writeclk_inv),
    
    .EXT_18K                (1'b0),
    .FIFO_EN                (1'b1),
    .PEEK_MODE              (peek),
    .PORTA_PROG             (8'b11110000),
    .PORTB_PROG             (8'b00001111),
    .WIDTH_EXT_MODE23       (1'b0),
    .WIDTH_EXT_MODE01       (1'b0)
)

u0_emb18k_core (
    .a_addr_ext             (),
    .b_addr_ext             (),
    
    .c1r4_aa                (),
    .c1r4_ab                (),
    .c1r4_cea               (),
    .c1r4_ceb               (),
    .c1r4_clka              (),
    .c1r4_clkb              (),
    .c1r4_da                (),
    .c1r4_db                (),
    .c1r4_rstna             (),
    .c1r4_rstnb             (),
    .c1r4_wea               (),
    .c1r4_web               (),
    .c1r4_user_ena          (),
    .c1r4_user_enb          (),
    
    .c1r3_aa                (),
    .c1r3_ab                (),
    .c1r3_cea               (),
    .c1r3_ceb               (),
    .c1r3_clka              (),
    .c1r3_clkb              (),
    .c1r3_da                (),
    .c1r3_db                (),
    .c1r3_rstna             (),
    .c1r3_rstnb             (),
    .c1r3_wea               (),
    .c1r3_web               (),
    .c1r3_user_ena          (),
    .c1r3_user_enb          (),
    
    .c1r2_aa                (),
    .c1r2_ab                (),
    .c1r2_cea               (),
    .c1r2_ceb               (),
    .c1r2_clka              (),
    .c1r2_clkb              (),
    .c1r2_da                (),
    .c1r2_db                (),
    .c1r2_rstna             (),
    .c1r2_rstnb             (),
    .c1r2_wea               (),
    .c1r2_web               (),
    .c1r2_user_ena          (),
    .c1r2_user_enb          (),    
    
    .c1r1_aa                (),
    .c1r1_ab                (),
    .c1r1_cea               (),
    .c1r1_ceb               (),
    .c1r1_clka              (readclk),
    .c1r1_clkb              (writeclk),
    .c1r1_da                (),
    .c1r1_db                (datain),
    .c1r1_rstna             (reset),
    .c1r1_rstnb             (1'b1),
    .c1r1_wea               (),
    .c1r1_web               (),
    .c1r1_user_ena          (regce),
    .c1r1_user_enb          (regce),
    
    .rd_mem_n               (rd_mem_n),
    .rptr                   (rptr[13:0]),
    .wptr                   (wptr[13:0]),
    .wr_mem_n               (wr_mem_n),      
    .peek_en                (peek_en),
    .peek_rd_en             (peek_rd_en),
    
    .c1r4_q                 (),
    .c1r3_q                 (),
    .c1r2_q                 (),
    .c1r1_q                 (dataout),
    .eccindberr             (1'b0),
    .eccinsberr             (1'b0),
    .eccoutdberr            (),
    .eccoutsberr            (),
    .err_addr               () 
);    
    
endmodule // FIFO5K

// end of FIFO5K 

module FIFO9K (dout, doutp, din, dinp, writeclk, readclk, writeen, readen, reset, regce, 
            writesave, writedrop, full, empty, almostfull, almostempty, overflow, underflow, writedropflag);

    output [31:0] dout;
    output [3:0] doutp;
    output full, empty;
    output almostfull, almostempty;
    output overflow, underflow;
    output writedropflag;
    
    input [31:0] din;
    input [3:0] dinp;
    input writeclk, readclk;
    input writeen, readen;
    input reset, regce;
    input writesave, writedrop;

    parameter almostemptyth = 13'b0;
    parameter almostfullth = 13'b0;
    parameter writewidth = 1;
    parameter readwidth = 1;
    parameter outreg = 0;
    parameter peek = 1'b0;
    parameter readclk_inv = 1'b0;
    parameter writeclk_inv = 1'b0;
    parameter use_parity = 0;
    
    reg finish_error = 0;
    
    initial begin
    
        if (peek == 1'b1 && outreg == 0) begin
            $display("DRC Error : outreg = 0 is invalid when peek is set to 1 on FIFO9K instance %m.");
            finish_error = 1;
        end
    
        case (readwidth)
            1: begin
                case (writewidth)
                    1, 2, 4, 9, 18: ;
                    default : begin
                        $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18.", readwidth);
                        finish_error = 1;
                    end
                endcase
            end
            
            2, 4, 18: begin
                case (writewidth)
                    1, 2, 4, 9, 18, 36: ;
                    default : begin
                        $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18, 36.", readwidth);
                        finish_error = 1;
                    end
                endcase
            end
            9: begin
                case (writewidth)
                    1, 2, 4, 36: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 9, 18.", readwidth);
                            finish_error = 1;
                        end
                    end
                    9, 18: ;
                    default : begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 9, 18.", readwidth);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18, 36.", readwidth);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            36: begin
                case (writewidth)
                    1: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 18, 36.", readwidth);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 2, 4, 9, 18, 36.", readwidth);
                            finish_error = 1;
                        end
                    end
                    2, 4, 9: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 18, 36.", readwidth);
                            finish_error = 1;
                        end
                    end
                    
                    18, 36: ;
                    default : begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 18, 36.", readwidth);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute writewidth are 2, 4, 9, 18, 36.", readwidth);
                            finish_error = 1;
                        end
                    end
                endcase
            end
    
            default: begin
                $display("Attribute Syntax Error : The attribute readwidth on FIFO9K instance %m is set to %d, Legal value for attribute readwidth are 1, 2, 4, 9, 18, 36.", readwidth);
                finish_error = 1;
            end
        endcase
        
        //if (finish_error == 1)
        //    $finish;
    end // end initial    
    
    parameter depth_extension = (readwidth == 36 || writewidth == 36) ? 1'b0 : 1'b1;
    parameter width_extension = (depth_extension == 1'b1) ? 1'b0 : 1'b1;

    parameter read_sel =    (readwidth == 1) ? 4'b1111 : 
                            (readwidth == 2) ? ((depth_extension == 1'b0) ? 4'b1111 : 4'b1110) :
                            (readwidth == 4) ? ((depth_extension == 1'b0) ? 4'b1110 : 4'b1100) :
                            (readwidth == 9) ? ((depth_extension == 1'b0) ? 4'b1100 : 4'b1000) :
                            (readwidth == 18) ? ((depth_extension == 1'b0) ? 4'b1000 : 4'b0000) :
                            (readwidth == 36) ? 4'b0000 : 4'bxxxx;
                           
    parameter write_sel =   (writewidth == 1) ? 4'b1111 : 
                            (writewidth == 2) ? ((depth_extension == 1'b0) ? 4'b1111 : 4'b1110) :
                            (writewidth == 4) ? ((depth_extension == 1'b0) ? 4'b1110 : 4'b1100) :
                            (writewidth == 9) ? ((depth_extension == 1'b0) ? 4'b1100 : 4'b1000) :
                            (writewidth == 18) ? ((depth_extension == 1'b0) ? 4'b1000 : 4'b0000) :                                
                            (writewidth == 36) ? 4'b0000 : 4'bxxxx;    

    parameter readwidth_5k =    (readwidth == 1) ? 1 : 
                                (readwidth == 2) ? ((depth_extension == 1'b0) ? 1 : 2) :
                                (readwidth == 4) ? ((depth_extension == 1'b0) ? 2 : 4) :
                                (readwidth == 9) ? ((depth_extension == 1'b0) ? 4 : 9) :
                                (readwidth == 18) ? ((depth_extension == 1'b0) ? 9 : 18) :
                                (readwidth == 36) ? 18 : 18;
                            
    parameter writewidth_5k =   (writewidth == 1) ? 1 : 
                                (writewidth == 2) ? ((depth_extension == 1'b0) ? 1 : 2) :
                                (writewidth == 4) ? ((depth_extension == 1'b0) ? 2 : 4) :
                                (writewidth == 9) ? ((depth_extension == 1'b0) ? 4 : 9) :
                                (writewidth == 18) ? ((depth_extension == 1'b0) ? 9 : 18) :
                                (writewidth == 36) ? 18 : 18;
                                
    parameter read_data_width_5k =  (readwidth_5k == 1) ? 1 : 
                                    (readwidth_5k == 2) ? 2 :
                                    (readwidth_5k == 4) ? 4 :
                                    (readwidth_5k == 9) ? 8 :
                                    (readwidth_5k == 18) ? 16 : 0;
                                
    parameter write_data_width_5k = (writewidth_5k == 1) ? 1 : 
                                    (writewidth_5k == 2) ? 2 :
                                    (writewidth_5k == 4) ? 4 :
                                    (writewidth_5k == 9) ? 8 :
                                    (writewidth_5k == 18) ? 16 : 0;

    parameter prog_full = (almostfullth + peek * 2) * write_data_width_5k;
    parameter prog_empty = (almostemptyth - peek * 2) * read_data_width_5k;                                    

    parameter EXT_18K = 1'b0;
                                
    wire rd_mem_n;
    wire [13:0]	rptr;
    wire [13:0]	wptr;
    wire wr_mem_n;

    wire peek_en;
    wire peek_rd_en;

/*    wire [17:0] datain_bnk1 =   (writewidth_5k == 18) ? {dinp[1:0], din[15:0]} : 
                                (writewidth_5k == 9) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                                (writewidth_5k == 4) ? {1'bx, 1'bx, {4{din[3:0]}}} :
                                (writewidth_5k == 2) ? {1'bx, 1'bx, {8{din[1:0]}}} :
                                (writewidth_5k == 1) ? {1'bx, 1'bx, {16{din[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;
    
    wire [17:0] datain_bnk2 =   (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx: {dinp[3:2], din[31:16]}) : 
                                (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {dinp[1], dinp[1], din[15:8], din[15:8]}) :
                                (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{din[7:4]}}}) :
                                (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx: {1'bx, 1'bx, {8{din[3:2]}}}) :
                                (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
*////
    wire [17:0] datain_bnk1 = (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? {dinp[1:0], din[15:0]}:
                                                      (writewidth_5k <= readwidth_5k) ? {dinp[1:0], din[15:0]}:
                                                      (readwidth_5k == 1) ? {dinp[2],dinp[0],din[30], din[28], din[26], din[24], din[22], din[20], din[18], din[16],din[14], din[12], din[10], din[8], din[6], din[4], din[2], din[0]}:
                                                      (readwidth_5k == 2) ? {dinp[2],dinp[0],din[29:28],din[25:24],din[21:20],din[17:16],din[13:12],din[9:8],din[5:4],din[1:0]}:
                                                      (readwidth_5k == 4) ? {dinp[2],dinp[0],din[27:24],din[19:16],din[11:8],din[3:0]}:
                                                      (readwidth_5k == 9) ? {dinp[2],dinp[0], din[23:16], din[7:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                                                      (writewidth_5k <= readwidth_5k) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                                                      (readwidth_5k == 1) ? {dinp[0],dinp[0],din[14], din[12], din[10], din[8], din[6], din[4], din[2], din[0],din[14], din[12], din[10], din[8], din[6], din[4], din[2], din[0]}:
                                                      (readwidth_5k == 2) ? {dinp[0],dinp[0],din[13:12],din[9:8],din[5:4],din[1:0],din[13:12],din[9:8],din[5:4],din[1:0]}:
                                                      (readwidth_5k == 4) ? {dinp[0],dinp[0],din[11:8],din[3:0],din[11:8],din[3:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (writewidth_5k == 4) ? {1'bx, 1'bx, {4{din[3:0]}}} :
                               (writewidth_5k == 2) ? {1'bx, 1'bx, {8{din[1:0]}}} :
                               (writewidth_5k == 1) ? {1'bx, 1'bx, {16{din[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;

    wire [17:0] datain_bnk2 = (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[3:2], din[31:16]}:
                                                      (readwidth_5k == 1) ? {dinp[3],dinp[1],din[31], din[29], din[27], din[25], din[23], din[21], din[19], din[17],din[15], din[13], din[11], din[9], din[7], din[5], din[3], din[1]}:
                                                      (readwidth_5k == 2) ? {dinp[3],dinp[1],din[31:30],din[27:26],din[23:22],din[19:18],din[15:14],din[11:10],din[7:6],din[3:2]}:
                                                      (readwidth_5k == 4) ? {dinp[3],dinp[1],din[31:28],din[23:20],din[15:12],din[7:4]}:
                                                      (readwidth_5k == 9) ? {dinp[3],dinp[1], din[31:24], din[15:8]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[1], dinp[1], din[15:8], din[15:8]} :
                                                      (readwidth_5k == 1) ? {dinp[1],dinp[1],din[15], din[13], din[11], din[9], din[7], din[5], din[3], din[1],din[15], din[13], din[11], din[9], din[7], din[5], din[3], din[1]}:
                                                      (readwidth_5k == 2) ? {dinp[1],dinp[1],din[15:14],din[11:10],din[7:6],din[3:2],din[15:14],din[11:10],din[7:6],din[3:2]}:
                                                      (readwidth_5k == 4) ? {dinp[1],dinp[1],din[15:12],din[7:4],din[15:12],din[7:4]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{din[7:4]}}}) :
                               (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[3:2]}}}) :
                               (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;							
								
/*								
    wire [17:0] dataout_bnk1;
    wire [17:0] dataout_bnk2;

    assign doutp[3] = (depth_extension == 1'b1) ?   1'bx : dataout_bnk2[17];
    assign doutp[1] = (depth_extension == 1'b1) ?   ((readwidth_5k == 18) ? dataout_bnk1[17] : 
                                                                            dataout_bnk2[8]) :
                                                    (readwidth_5k == 18) ?  dataout_bnk1[17] : 
                                                                            1'bx;
    assign doutp[2] = (depth_extension == 1'b1) ?   1'bx : 
                                                    ((readwidth_5k == 18) ? dataout_bnk2[16] : 
                                                                            dataout_bnk2[8]);
    assign doutp[0] = (readwidth_5k == 18) ? dataout_bnk1[16] : dataout_bnk1[8];    

    assign dout[7:0] = dataout_bnk1[7:0];
    assign dout[15:8] =  (readwidth_5k == 18) ? dataout_bnk1[15:8] : 
                        (depth_extension == 1'b1) ? 8'bxxxxxxxx : 
                                                    dataout_bnk2[7:0];
    assign dout[31:16] = (readwidth_5k == 18 && depth_extension == 1'b0) ? dataout_bnk2[15:0] : 16'bxxxxxxxxxxxxxxxx;
*/////

    wire [17:0] dataout_bnk1;
    wire [17:0] dataout_bnk2;
	
    assign doutp[3] = (depth_extension == 1'b1) ? 1'bx : dataout_bnk2[17];
    assign doutp[1] = (depth_extension == 1'b1) ? dataout_bnk1[17] :((readwidth_5k == 9) ? dataout_bnk2[8] :((readwidth_5k == 18) ? ((writewidth_5k == 18) ?dataout_bnk1[17]: dataout_bnk2[16]) : dataout_bnk2[8]));
    assign doutp[2] = (depth_extension == 1'b1) ? 1'bx : ((readwidth_5k == writewidth_5k) ? dataout_bnk2[16]:dataout_bnk1[17]);
    assign doutp[0] = (readwidth_5k == 18) ? dataout_bnk1[16] : dataout_bnk1[8];

    assign dout = readwidth_5k==1 ? {30'h0,dataout_bnk2[0],dataout_bnk1[0]} :
                  readwidth_5k==2 ? {28'h0,dataout_bnk2[1:0],dataout_bnk1[1:0]} :
                  readwidth_5k==4 ? {24'h0,dataout_bnk2[3:0],dataout_bnk1[3:0]} :
                  readwidth_5k==9 ? ((depth_extension == 1'b1) ? {16'h0,dataout_bnk2[7:0],dataout_bnk1[7:0]} :
                                   (writewidth_5k >= readwidth_5k) ?{16'h0,dataout_bnk2[7:0],dataout_bnk1[7:0]} :                            
                                   (writewidth_5k == 4) ? {dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (writewidth_5k == 2) ? {dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (writewidth_5k == 1) ? {dataout_bnk2[7],dataout_bnk1[7],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk2[0],dataout_bnk1[0]}:{dataout_bnk2[15:0],dataout_bnk1[15:0]  }) :
                 
                  readwidth_5k==18 ? ((depth_extension == 1'b1) ? {dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (writewidth_5k >= readwidth_5k) ?{dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (writewidth_5k == 9) ? {dataout_bnk2[15:8],dataout_bnk1[15:8],dataout_bnk2[7:0],dataout_bnk1[7:0]  }:
                                   (writewidth_5k == 4) ? {dataout_bnk2[15:12],dataout_bnk1[15:12],dataout_bnk2[11:8],dataout_bnk1[11:8],dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (writewidth_5k == 2) ? {dataout_bnk2[15:14],dataout_bnk1[15:14],dataout_bnk2[13:12],dataout_bnk1[13:12],dataout_bnk2[11:10],dataout_bnk1[11:10],dataout_bnk2[9:8],dataout_bnk1[9:8],dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (writewidth_5k == 1) ? {dataout_bnk2[15],dataout_bnk1[15],dataout_bnk2[14],dataout_bnk1[14],dataout_bnk2[13],dataout_bnk1[13],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk2[9],dataout_bnk1[9],dataout_bnk2[8],dataout_bnk1[8],dataout_bnk2[7],dataout_bnk1[7],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk2[0],dataout_bnk1[0]}:{dataout_bnk2[15:0],dataout_bnk1[15:0]  }) :
                 32'hxxxx_xxxx; 
FIFOCTRL18KV1 # (
	.USR_PF		({1'b0, prog_full}),
	.USR_PE		({1'b0, prog_empty}),
	.PEEK_MODE	(peek),
	.FIFO_EN	(1'b1),
	.R_WIDTH	(read_sel),
	.W_WIDTH	(write_sel),
	.DEPTH_EXT_MODE	({EXT_18K, depth_extension})
)
u0_fifo_ctrl (
	.rst_n		(reset),
	.rd_req_n	(readen),
	.wr_req_n	(writeen),
	.clka		(readclk),
	.clkb		(writeclk),
	.write_drop	(writedrop),
	.write_save	(writesave),


	.full		(full),
	.empty		(empty),
	.prog_full	(almostfull),
	.prog_empty	(almostempty),
	.wptr		(wptr[13:0]),
	.rptr		(rptr[13:0]),
	.wr_mem_n	(wr_mem_n),
	.rd_mem_n	(rd_mem_n),
	.overflow	(overflow),
	.underflow	(underflow),
    .wrdp_rd_flag(writedropflag),
	.peek_en	(peek_en),
    .peek_rd_en (peek_rd_en)    
);

BRAM18KV1 # (
    .DEPTH_EXT_MODE23       (1'b0),
    .DEPTH_EXT_MODE01       (depth_extension),
    .ECC_DEC_EN             (1'b0),
    .ECC_ENC_EN             (1'b0),
    
    .EMB5K_4_MODEA_SEL      (),
    .EMB5K_4_MODEB_SEL      (),
    .EMB5K_4_PORTA_BYPASS   (),
    .EMB5K_4_PORTA_CE       (),
    .EMB5K_4_PORTA_REG_OUT  (),
    .EMB5K_4_PORTA_WR_MODE  (),
    .EMB5K_4_PORTA_CKINV    (),
    .EMB5K_4_PORTB_BYPASS   (),
    .EMB5K_4_PORTB_CE       (),
    .EMB5K_4_PORTB_REG_OUT  (),
    .EMB5K_4_PORTB_WR_MODE  (),
    .EMB5K_4_PORTB_CKINV    (),
    
    .EMB5K_3_MODEA_SEL      (),
    .EMB5K_3_MODEB_SEL      (),
    .EMB5K_3_PORTA_BYPASS   (),
    .EMB5K_3_PORTA_CE       (),
    .EMB5K_3_PORTA_REG_OUT  (),
    .EMB5K_3_PORTA_WR_MODE  (),
    .EMB5K_3_PORTA_CKINV    (),
    .EMB5K_3_PORTB_BYPASS   (),
    .EMB5K_3_PORTB_CE       (),
    .EMB5K_3_PORTB_REG_OUT  (),
    .EMB5K_3_PORTB_WR_MODE  (),
    .EMB5K_3_PORTB_CKINV    (),
    
    .EMB5K_2_MODEA_SEL      (read_sel),
    .EMB5K_2_MODEB_SEL      (write_sel),
    .EMB5K_2_PORTA_BYPASS   (1'b0),
    .EMB5K_2_PORTA_CE       (1'b1),
    .EMB5K_2_PORTA_REG_OUT  (outreg),
    .EMB5K_2_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_2_PORTA_CKINV    (readclk_inv),
    .EMB5K_2_PORTB_BYPASS   (1'b0),
    .EMB5K_2_PORTB_CE       (1'b1),
    .EMB5K_2_PORTB_REG_OUT  (),
    .EMB5K_2_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_2_PORTB_CKINV    (writeclk_inv),
    
    .EMB5K_1_MODEA_SEL      (read_sel),
    .EMB5K_1_MODEB_SEL      (write_sel),
    .EMB5K_1_PORTA_BYPASS   (1'b0),
    .EMB5K_1_PORTA_CE       (1'b1),
    .EMB5K_1_PORTA_REG_OUT  (outreg),
    .EMB5K_1_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_1_PORTA_CKINV    (readclk_inv),
    .EMB5K_1_PORTB_BYPASS   (1'b0),
    .EMB5K_1_PORTB_CE       (1'b1),
    .EMB5K_1_PORTB_REG_OUT  (),
    .EMB5K_1_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_1_PORTB_CKINV    (writeclk_inv),  

    .EXT_18K                (EXT_18K),
    .FIFO_EN                (1'b1),
    .PEEK_MODE              (peek),
    .PORTA_PROG             (8'b11110000),
    .PORTB_PROG             (8'b00001111),
    .WIDTH_EXT_MODE23       (1'b0),
    .WIDTH_EXT_MODE01       (width_extension)
)
u0_emb18k_core ( 
    .a_addr_ext             (),
    .b_addr_ext             (),
    
    .c1r4_aa                (),
    .c1r4_ab                (),
    .c1r4_cea               (),
    .c1r4_ceb               (),
    .c1r4_clka              (),
    .c1r4_clkb              (),
    .c1r4_da                (),
    .c1r4_db                (),
    .c1r4_rstna             (),
    .c1r4_rstnb             (),
    .c1r4_wea               (),
    .c1r4_web               (),
    .c1r4_user_ena          (),
    .c1r4_user_enb          (),
    
    .c1r3_aa                (),
    .c1r3_ab                (),
    .c1r3_cea               (),
    .c1r3_ceb               (),
    .c1r3_clka              (),
    .c1r3_clkb              (),
    .c1r3_da                (),
    .c1r3_db                (),
    .c1r3_rstna             (),
    .c1r3_rstnb             (),
    .c1r3_wea               (),
    .c1r3_web               (),
    .c1r3_user_ena          (),
    .c1r3_user_enb          (),
    
    .c1r2_aa                (),
    .c1r2_ab                (),
    .c1r2_cea               (),
    .c1r2_ceb               (),
    .c1r2_clka              (readclk),
    .c1r2_clkb              (writeclk),
    .c1r2_da                (),
    .c1r2_db                (datain_bnk2),
    .c1r2_rstna             (1'b1),
    .c1r2_rstnb             (1'b1),
    .c1r2_wea               (),
    .c1r2_web               (),
    .c1r2_user_ena          (regce),
    .c1r2_user_enb          (regce),    
    
    .c1r1_aa                (),
    .c1r1_ab                (),
    .c1r1_cea               (),
    .c1r1_ceb               (),
    .c1r1_clka              (readclk),
    .c1r1_clkb              (writeclk),
    .c1r1_da                (),
    .c1r1_db                (datain_bnk1),
    .c1r1_rstna             (reset),
    .c1r1_rstnb             (1'b1),
    .c1r1_wea               (),
    .c1r1_web               (),
    .c1r1_user_ena          (regce),
    .c1r1_user_enb          (regce),
    
    .rd_mem_n               (rd_mem_n),
    .rptr                   (rptr[13:0]),
    .wptr                   (wptr[13:0]),
    .wr_mem_n               (wr_mem_n),      
    .peek_en                (peek_en),
    .peek_rd_en             (peek_rd_en),
    
    .c1r4_q                 (),
    .c1r3_q                 (),
    .c1r2_q                 (dataout_bnk2),
    .c1r1_q                 (dataout_bnk1),
    .eccindberr             (1'b0),
    .eccinsberr             (1'b0),
    .eccoutdberr            (),
    .eccoutsberr            (),
    .err_addr               () 
);    
    
endmodule // FIFO9K

// end of FIFO9K 

module FIFO18K (dout, doutp, din, dinp, writeclk, readclk, writeen, readen, reset, regce, 
            writesave, writedrop, full, empty, almostfull, almostempty, overflow, underflow, 
            eccoutdberr, eccoutsberr, eccreadaddr, eccindberr, eccinsberr, writedropflag);

    output [63:0] dout;
    output [7:0] doutp;
    output full, empty;
    output almostfull, almostempty;
    output overflow, underflow;
    output eccoutdberr, eccoutsberr;
    output [7:0] eccreadaddr;
    output writedropflag;
    
    input [63:0] din;
    input [7:0] dinp;
    input writeclk, readclk;
    input writeen, readen;
    input reset, regce;
    input eccindberr, eccinsberr;
    input writesave, writedrop;

    parameter eccreaden = 0;
    parameter eccwriteen = 0;
    parameter almostemptyth = 14'b0;
    parameter almostfullth = 14'b0;
    parameter writewidth = 1;
    parameter readwidth = 1;
    parameter outreg = 0;
    parameter peek = 1'b0;
    parameter readclk_inv = 1'b0;
    parameter writeclk_inv = 1'b0;
    parameter use_parity = 0;
    
    reg finish_error = 0;
    
    initial begin
    
        if (peek == 1'b1 && outreg == 0) begin
            $display("DRC Error : outreg = 0 is invalid when peek is set to 1 on FIFO18K instance %m.");
            finish_error = 1;
        end
    
        case (readwidth)
            1: begin
                case (writewidth)
                    1, 2, 4, 9, 18: ;
                    default : begin
                        $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18.", readwidth);
                        finish_error = 1;
                    end
                endcase
            end
            
            2: begin
                case (writewidth)
                    1, 2, 4, 9, 18: ;
                    default : begin
                        $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18.", readwidth);
                        finish_error = 1;
                    end
                endcase
            end
            
            4: begin
                case (writewidth)
                    1, 2, 4, 9, 18, 36, 72: ;
                    default : begin
                        $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18, 36, 72.", readwidth);
                        finish_error = 1;
                    end
                endcase
            end
            9, 18: begin
                case (writewidth)
                    1, 2, 4, 36, 72: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 9, 18.", readwidth);
                            finish_error = 1;
                        end
                    end
                    9, 18: ;
                    default : begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 9, 18.", readwidth);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 1, 2, 4, 9, 18, 36, 72.", readwidth);
                            finish_error = 1;
                        end
                    end
                endcase
            end
            36, 72: begin
                case (writewidth)
                    1, 2: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 36, 72.", readwidth);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 4, 9, 18, 36, 72.", readwidth);
                            finish_error = 1;
                        end
                    end
                    4, 9, 18: begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 36, 72.", readwidth);
                            finish_error = 1;
                        end
                    end
                    
                    36, 72: ;
                    default : begin
                        if (use_parity == 1) begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 36, 72.", readwidth);
                            finish_error = 1;
                        end
                        else begin
                            $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute writewidth are 4, 9, 18, 36, 72.", readwidth);
                            finish_error = 1;
                        end
                    end
                endcase
            end
    
            default: begin
                $display("Attribute Syntax Error : The attribute readwidth on FIFO18K instance %m is set to %d, Legal value for attribute readwidth are 1, 2, 4, 9, 18, 36, 72.", readwidth);
                finish_error = 1;
            end
        endcase
        
        //if (finish_error == 1)
        //    $finish;
    end // end initial
        
    parameter depth_extension = (readwidth == 72 || readwidth == 36 
                                || writewidth == 72 || writewidth == 36) ? 1'b0 : 1'b1;
    parameter width_extension = (depth_extension == 1'b1) ? 1'b0 : 1'b1;
    
    parameter readwidth_5k =    (readwidth == 1) ? 1 : 
                                (readwidth == 2) ? 2 :
                                (readwidth == 4) ? ((depth_extension == 1'b0) ? 1 : 4) :
                                (readwidth == 9) ? ((depth_extension == 1'b0) ? 2 : 9) :
                                (readwidth == 18) ? ((depth_extension == 1'b0) ? 4 : 18) :
                                (readwidth == 36) ? 9 :
                                (readwidth == 72) ? 18 : 18;
                            
    parameter writewidth_5k =   (writewidth == 1) ? 1 : 
                                (writewidth == 2) ? 2 :
                                (writewidth == 4) ? ((depth_extension == 1'b0) ? 1 : 4) :
                                (writewidth == 9) ? ((depth_extension == 1'b0) ? 2 : 9) :
                                (writewidth == 18) ? ((depth_extension == 1'b0) ? 4 : 18) :
                                (writewidth == 36) ? 9 :
                                (writewidth == 72) ? 18 : 18;

    parameter read_sel =    (readwidth_5k == 1) ? 4'b1111 : 
                            (readwidth_5k == 2) ? 4'b1110 :
                            (readwidth_5k == 4) ? 4'b1100 :
                            (readwidth_5k == 9) ? 4'b1000 :
                            (readwidth_5k == 18) ? 4'b0000 : 4'bxxxx;
                           
    parameter write_sel =   (writewidth_5k == 1) ? 4'b1111 : 
                            (writewidth_5k == 2) ? 4'b1110 :
                            (writewidth_5k == 4) ? 4'b1100 :
                            (writewidth_5k == 9) ? 4'b1000 :
                            (writewidth_5k == 18) ? 4'b0000 : 4'bxxxx;
                            
    parameter read_data_width_5k =  (readwidth_5k == 1) ? 1 : 
                                    (readwidth_5k == 2) ? 2 :
                                    (readwidth_5k == 4) ? 4 :
                                    (readwidth_5k == 9) ? 8 :
                                    (readwidth_5k == 18) ? 16 : 0;
                                
    parameter write_data_width_5k = (writewidth_5k == 1) ? 1 : 
                                    (writewidth_5k == 2) ? 2 :
                                    (writewidth_5k == 4) ? 4 :
                                    (writewidth_5k == 9) ? 8 :
                                    (writewidth_5k == 18) ? 16 : 0;

    parameter prog_full = (almostfullth + peek * 2) * write_data_width_5k;
    parameter prog_empty = (almostemptyth - peek * 2) * read_data_width_5k; 
                            
    parameter ext_18k = 1'b1;
                
    wire rd_mem_n;
    wire [13:0]	rptr;
    wire [13:0]	wptr;
    wire wr_mem_n;

    wire peek_en;
    wire peek_rd_en;

 /*   wire [17:0] datain_bnk1 =   (writewidth_5k == 18) ? {dinp[1:0], din[15:0]} : 
                                (writewidth_5k == 9) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                                (writewidth_5k == 4) ? {1'bx, 1'bx, {4{din[3:0]}}} :
                                (writewidth_5k == 2) ? {1'bx, 1'bx, {8{din[1:0]}}} :
                                (writewidth_5k == 1) ? {1'bx, 1'bx, {16{din[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;
    
    wire [17:0] datain_bnk2 =   (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {dinp[3:2], din[31:16]}) : 
                                (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {dinp[1], dinp[1], din[15:8], din[15:8]}) :
                                (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{din[7:4]}}}) :
                                (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[3:2]}}}) :
                                (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;

    wire [17:0] datain_bnk3 =   (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx :  {dinp[5:4], din[47:32]}) : 
                                (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {dinp[2], dinp[2], din[23:16], din[23:16]}) :
                                (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{din[11:8]}}}) :
                                (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[5:4]}}}) :
                                (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[2]}}}) : 18'bxxxxxxxxxxxxxxxxxx;

    wire [17:0] datain_bnk4 =   (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {dinp[7:6], din[63:48]}) : 
                                (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {dinp[3], dinp[3], din[31:24], din[31:24]}) :
                                (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {4{din[15:12]}}}) :
                                (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[7:6]}}}) :
                                (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[3]}}}) : 18'bxxxxxxxxxxxxxxxxxx;                                
                                
    wire [17:0] dataout_bnk1;
    wire [17:0] dataout_bnk2;
    wire [17:0] dataout_bnk3;
    wire [17:0] dataout_bnk4;
    
    assign doutp[7:4] = (depth_extension == 1'b1) ? 4'bxxxx : 
                        (readwidth_5k == 18) ? {dataout_bnk4[17], dataout_bnk4[16], dataout_bnk3[17], dataout_bnk3[16]} :
                        4'bxxxx;

    assign doutp[3:2] = (depth_extension == 1'b1) ? 2'bxx : 
                        (readwidth_5k == 18) ?  {dataout_bnk2[17], dataout_bnk2[16]} : 
                                                {dataout_bnk4[8], dataout_bnk3[8]};

    assign doutp[1:0] = (depth_extension == 1'b1) ? ((readwidth_5k == 18) ? {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                                            {1'bx, dataout_bnk1[8]}) : 
                        (readwidth_5k == 18) ?    {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                {dataout_bnk2[8], dataout_bnk1[8]};

    assign dout[63:32] =    (depth_extension == 1'b1) ? 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx : 
                            (readwidth_5k == 18) ? {dataout_bnk4[15:0], dataout_bnk3[15:0]} :
                            32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;

    assign dout[31:16] =    (depth_extension == 1'b1) ? 16'bxxxxxxxxxxxxxxxx : 
                            (readwidth_5k == 18) ?    dataout_bnk2[15:0] : 
                                                    {dataout_bnk4[7:0], dataout_bnk3[7:0]};                        

    assign dout[15:8] =     (depth_extension == 1'b1) ? ((readwidth_5k == 18) ? dataout_bnk1[15:8] : 
                                                                                8'bxxxxxxxx) : 
                            (readwidth_5k == 18) ?  dataout_bnk1[15:8] : 
                                                    dataout_bnk2[7:0];
                                                
    assign dout[7:0] =      dataout_bnk1[7:0]; 
 */
    wire [17:0] datain_bnk1 = (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? {dinp[1:0], din[15:0]}:
                                                      (writewidth_5k <= readwidth_5k) ? {dinp[1:0], din[15:0]}:
                                                      (readwidth_5k == 1) ? {dinp[4],dinp[0],din[60], din[56], din[52], din[48], din[44], din[40], din[36], din[32],din[28], din[24], din[20], din[16], din[12], din[8], din[4], din[0]}:
                                                      (readwidth_5k == 2) ? {dinp[4],dinp[0],din[57:56],din[49:48],din[41:40],din[33:32],din[25:24],din[17:16],din[9:8],din[1:0]}:
                                                      (readwidth_5k == 4) ? {dinp[4],dinp[0],din[51:48],din[35:32],din[19:16],din[3:0]}:
                                                      (readwidth_5k == 9) ? {dinp[4],dinp[0], din[39:32], din[7:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                                                      (writewidth_5k <= readwidth_5k) ? {dinp[0], dinp[0], din[7:0], din[7:0]} :
                                                      (readwidth_5k == 1) ? {dinp[0],dinp[0],din[28], din[24], din[20], din[16], din[12], din[8], din[4], din[0],din[28], din[24], din[20], din[16], din[12], din[8], din[4], din[0]}:
                                                      (readwidth_5k == 2) ? {dinp[0],dinp[0],din[25:24],din[17:16],din[9:8],din[1:0],din[25:24],din[17:16],din[9:8],din[1:0]}:
                                                      (readwidth_5k == 4) ? {dinp[0],dinp[0],din[19:16],din[3:0],din[19:16],din[3:0]}:18'bxxxxxxxxxxxxxxxxxx): 
                               (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? {1'bx, 1'bx, {4{din[3:0]}}} :
							                          (writewidth_5k <= readwidth_5k) ? {1'bx, 1'bx, {4{din[3:0]}}} :
                                                      (readwidth_5k == 1) ? {1'bx, 1'bx, {4{din[12], din[8], din[4], din[0]}}}:
                                                      (readwidth_5k == 2) ? {1'bx, 1'bx, {4{din[9:8],din[1:0]}}} :18'bxxxxxxxxxxxxxxxxxx): 
                                                      
                               (writewidth_5k == 2) ? {1'bx, 1'bx, {8{din[1:0]}}} :
                               (writewidth_5k == 1) ? {1'bx, 1'bx, {16{din[0]}}} : 18'bxxxxxxxxxxxxxxxxxx;


    wire [17:0] datain_bnk2 = (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[3:2], din[31:16]}:
                                                      (readwidth_5k == 1) ? {dinp[5],dinp[1],din[61], din[57], din[53], din[49], din[45], din[41], din[37], din[33],din[29], din[25], din[21], din[17], din[13], din[9], din[5], din[1]}:
                                                      (readwidth_5k == 2) ? {dinp[5],dinp[1],din[59:58],din[51:50],din[43:42],din[35:34],din[27:26],din[19:18],din[11:10],din[3:2]}:
                                                      (readwidth_5k == 4) ? {dinp[5],dinp[1],din[55:52],din[39:36],din[23:20],din[7:4]}:
                                                      (readwidth_5k == 9) ? {dinp[5],dinp[1], din[47:40], din[15:8]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[1], dinp[1], din[15:8], din[15:8]} :
                                                      (readwidth_5k == 1) ? {dinp[1],dinp[1],din[29], din[25], din[21], din[17], din[13], din[9], din[5], din[1],din[29], din[25], din[21], din[17], din[13], din[9], din[5], din[1]}:
                                                      (readwidth_5k == 2) ? {dinp[1],dinp[1],din[27:26],din[19:18],din[11:10],din[3:2],din[27:26],din[19:18],din[11:10],din[3:2]}:
                                                      (readwidth_5k == 4) ? {dinp[1],dinp[1],din[23:20],din[7:4],din[23:20],din[7:4]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {1'bx, 1'bx, {4{din[7:4]}}}: 
							                          (readwidth_5k == 1) ? {1'bx, 1'bx,{4{din[13], din[9], din[5], din[1]}}}:
                                                      (readwidth_5k == 2) ? {1'bx, 1'bx,{4{din[11:10],din[3:2]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[3:2]}}}) :
                               (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[1]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                        
						
   wire [17:0] datain_bnk3 = (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[5:4], din[47:32]}:
                                                      (readwidth_5k == 1) ? {dinp[6],dinp[2],din[62], din[58], din[54], din[50], din[46], din[42], din[38], din[34],din[30], din[26], din[22], din[18], din[14], din[10], din[6], din[2]}:
                                                      (readwidth_5k == 2) ? {dinp[6],dinp[2],din[61:60],din[53:52],din[45:44],din[37:36],din[29:28],din[21:20],din[13:12],din[5:4]}:
                                                      (readwidth_5k == 4) ? {dinp[6],dinp[2],din[59:56],din[43:40],din[27:24],din[11:8]}:
                                                      (readwidth_5k == 9) ? {dinp[6],dinp[2], din[55:48], din[23:16]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[2], dinp[2], din[23:16], din[23:16]} :
                                                      (readwidth_5k == 1) ? {dinp[2],dinp[2],din[30], din[26], din[22], din[18], din[14], din[10], din[6], din[2],din[30], din[26], din[22], din[18], din[14], din[10], din[6], din[2]}:
                                                      (readwidth_5k == 2) ? {dinp[2],dinp[2],din[29:28],din[21:20],din[13:12],din[5:4],din[29:28],din[21:20],din[13:12],din[5:4]}:
                                                      (readwidth_5k == 4) ? {dinp[2],dinp[2],din[27:24],din[11:8],din[27:24],din[11:8]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {1'bx, 1'bx, {4{din[11:8]}}} :
							                          (readwidth_5k == 1) ? {1'bx, 1'bx, {4{din[14], din[10], din[6], din[2]}}}:
                                                      (readwidth_5k == 2) ? {1'bx, 1'bx, {4{din[13:12],din[5:4]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[5:4]}}}) :
                               (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[2]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
                            
   wire [17:0] datain_bnk4 = (writewidth_5k == 18) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[7:6], din[63:48]}:
                                                      (readwidth_5k == 1) ? {dinp[7],dinp[3],din[63], din[59], din[55], din[51], din[47], din[43], din[39], din[35],din[31], din[27], din[23], din[19], din[15], din[11], din[7], din[3]}:
                                                      (readwidth_5k == 2) ? {dinp[7],dinp[3],din[63:62],din[55:54],din[47:46],din[39:38],din[31:30],din[23:22],din[15:14],din[7:6]}:
                                                      (readwidth_5k == 4) ? {dinp[7],dinp[3],din[63:60],din[47:44],din[31:28],din[15:12]}:
                                                      (readwidth_5k == 9) ? {dinp[7],dinp[3], din[63:56], din[31:24]}:18'bxxxxxxxxxxxxxxxxxx) : 
                               (writewidth_5k == 9) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {dinp[3], dinp[3], din[31:24], din[31:24]} :
                                                      (readwidth_5k == 1) ? {dinp[3],dinp[3],din[31], din[27], din[23], din[19], din[15], din[11], din[7], din[3],din[31], din[27], din[23], din[19], din[15], din[11], din[7], din[3]}:
                                                      (readwidth_5k == 2) ? {dinp[3],dinp[3],din[31:30],din[23:22],din[15:14],din[7:6],din[31:30],din[23:22],din[15:14],din[7:6]}:
                                                      (readwidth_5k == 4) ? {dinp[3],dinp[3],din[31:28],din[15:12],din[31:28],din[15:12]}:18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 4) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : (writewidth_5k <= readwidth_5k) ? {1'bx, 1'bx, {4{din[15:12]}}} :
							                          (readwidth_5k == 1) ? {1'bx, 1'bx, {4{din[15], din[11], din[7], din[3]}}}:
                                                      (readwidth_5k == 2) ? {1'bx, 1'bx, {4{din[15:14],din[7:6]}}}: 18'bxxxxxxxxxxxxxxxxxx) :
                               (writewidth_5k == 2) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {8{din[7:6]}}}) :
                               (writewidth_5k == 1) ? ((depth_extension == 1'b1) ? 18'bxxxxxxxxxxxxxxxxxx : {1'bx, 1'bx, {16{din[3]}}}) : 18'bxxxxxxxxxxxxxxxxxx;
 
 
    wire [7:0] doutp_buf0;
    wire [7:0] doutp_buf1;
	
    assign doutp = doutp_buf1;                      
    assign doutp_buf1 =  (depth_extension == 1'b1) ? doutp_buf0 :
                        (readwidth_5k <= writewidth_5k) ? doutp_buf0 :
                        (writewidth_5k == 9) ? {doutp_buf0[7], doutp_buf0[5], doutp_buf0[3], doutp_buf0[1], 
                                            doutp_buf0[6], doutp_buf0[4], doutp_buf0[2], doutp_buf0[0]} : doutp_buf0;
                                                                                                             
    wire [17:0] dataout_bnk1;
    wire [17:0] dataout_bnk2;
    wire [17:0] dataout_bnk3;
    wire [17:0] dataout_bnk4;
              
    assign doutp_buf0[7:4] = (depth_extension == 1'b1) ? 4'bxxxx : 
                            (depth_extension == 1'b1) ? 4'bxxxx : 
                            (readwidth_5k == 18) ?    {dataout_bnk4[17], dataout_bnk4[16], dataout_bnk3[17], dataout_bnk3[16]}
                                                    :4'bxxxx;

    assign doutp_buf0[3:2] = (depth_extension == 1'b1) ? 2'bxx : 
                            (depth_extension == 1'b1) ? ((readwidth_5k == 18) ? {dataout_bnk3[17], dataout_bnk3[16]} : 
                                                                                2'bxx) : 
                            (readwidth_5k == 18) ?    {dataout_bnk2[17], dataout_bnk2[16]} : 
                                                    {dataout_bnk4[8], dataout_bnk3[8]};

    assign doutp_buf0[1:0] = (depth_extension == 1'b1) ? ((readwidth_5k == 18) ? {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                                                {1'bx, dataout_bnk1[8]}) : 
                            (depth_extension == 1'b1) ? ((readwidth_5k == 18) ? {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                                                {dataout_bnk3[8], dataout_bnk1[8]}) : 
                            (readwidth_5k == 18) ?    {dataout_bnk1[17], dataout_bnk1[16]} : 
                                                    {dataout_bnk2[8], dataout_bnk1[8]};
                                                
	assign dout = readwidth_5k==1 ? {60'h0,dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]} :
                 readwidth_5k==2 ? {56'h0,dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]} :
                 readwidth_5k==4 ? ((depth_extension == 1'b1) ? {48'h0,dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]} :
				                   (writewidth_5k >= readwidth_5k) ? {48'h0,dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]} :                           
                                   (writewidth_5k == 2) ? {48'h0,dataout_bnk4[3:2],dataout_bnk3[3:2],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (writewidth_5k == 1) ? {48'h0,dataout_bnk4[3],dataout_bnk3[3],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk4[2],dataout_bnk3[2],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk4[1],dataout_bnk3[1],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]}: 
								   {48'h0,dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]}):
								   
                 readwidth_5k==9 ? ((depth_extension == 1'b1) ? {32'h0,dataout_bnk4[7:0],dataout_bnk3[7:0],dataout_bnk2[7:0],dataout_bnk1[7:0]} :
                                   (writewidth_5k >= readwidth_5k) ?{32'h0,dataout_bnk4[7:0],dataout_bnk3[7:0],dataout_bnk2[7:0],dataout_bnk1[7:0]} :                            
                                   (writewidth_5k == 4) ? {dataout_bnk4[7:4],dataout_bnk3[7:4],dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (writewidth_5k == 2) ? {dataout_bnk4[7:6],dataout_bnk3[7:6],dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk4[5:4],dataout_bnk3[5:4],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk4[3:2],dataout_bnk3[3:2],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (writewidth_5k == 1) ? {dataout_bnk4[7],dataout_bnk3[7],dataout_bnk2[7],dataout_bnk1[7],dataout_bnk4[6],dataout_bnk3[6],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk4[5],dataout_bnk3[5],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk4[4],dataout_bnk3[4],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk4[3],dataout_bnk3[3],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk4[2],dataout_bnk3[2],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk4[1],dataout_bnk3[1],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]}:
								   {dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0]  }) :
                 
                 readwidth_5k==18 ? ((depth_extension == 1'b1) ? {dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (writewidth_5k >= readwidth_5k) ?{dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0]  }:
                                   (writewidth_5k == 9) ? {dataout_bnk4[15:8],dataout_bnk3[15:8],dataout_bnk2[15:8],dataout_bnk1[15:8],dataout_bnk4[7:0],dataout_bnk3[7:0],dataout_bnk2[7:0],dataout_bnk1[7:0]  }:
                                   (writewidth_5k == 4) ? {dataout_bnk4[15:12],dataout_bnk3[15:12],dataout_bnk2[15:12],dataout_bnk1[15:12],dataout_bnk4[11:8],dataout_bnk3[11:8],dataout_bnk2[11:8],dataout_bnk1[11:8],dataout_bnk4[7:4],dataout_bnk3[7:4],dataout_bnk2[7:4],dataout_bnk1[7:4],dataout_bnk4[3:0],dataout_bnk3[3:0],dataout_bnk2[3:0],dataout_bnk1[3:0]  }:
                                   (writewidth_5k == 2) ? {dataout_bnk4[15:14],dataout_bnk3[15:14],dataout_bnk2[15:14],dataout_bnk1[15:14],dataout_bnk4[13:12],dataout_bnk3[13:12],dataout_bnk2[13:12],dataout_bnk1[13:12],dataout_bnk4[11:10],dataout_bnk3[11:10],dataout_bnk2[11:10],dataout_bnk1[11:10],dataout_bnk4[9:8],dataout_bnk3[9:8],dataout_bnk2[9:8],dataout_bnk1[9:8],dataout_bnk4[7:6],dataout_bnk3[7:6],dataout_bnk2[7:6],dataout_bnk1[7:6],dataout_bnk4[5:4],dataout_bnk3[5:4],dataout_bnk2[5:4],dataout_bnk1[5:4],dataout_bnk4[3:2],dataout_bnk3[3:2],dataout_bnk2[3:2],dataout_bnk1[3:2],dataout_bnk4[1:0],dataout_bnk3[1:0],dataout_bnk2[1:0],dataout_bnk1[1:0]  }:
                                   (writewidth_5k == 1) ? {dataout_bnk4[15],dataout_bnk3[15],dataout_bnk2[15],dataout_bnk1[15],dataout_bnk4[14],dataout_bnk3[14],dataout_bnk2[14],dataout_bnk1[14],dataout_bnk4[13],dataout_bnk3[13],dataout_bnk2[13],dataout_bnk1[13],dataout_bnk4[12],dataout_bnk3[12],dataout_bnk2[12],dataout_bnk1[12],dataout_bnk4[11],dataout_bnk3[11],dataout_bnk2[11],dataout_bnk1[11],dataout_bnk4[10],dataout_bnk3[10],dataout_bnk2[10],dataout_bnk1[10],dataout_bnk4[9],dataout_bnk3[9],dataout_bnk2[9],dataout_bnk1[9],dataout_bnk4[8],dataout_bnk3[8],dataout_bnk2[8],dataout_bnk1[8],dataout_bnk4[7],dataout_bnk3[7],dataout_bnk2[7],dataout_bnk1[7],dataout_bnk4[6],dataout_bnk3[6],dataout_bnk2[6],dataout_bnk1[6],dataout_bnk4[5],dataout_bnk3[5],dataout_bnk2[5],dataout_bnk1[5],dataout_bnk4[4],dataout_bnk3[4],dataout_bnk2[4],dataout_bnk1[4],dataout_bnk4[3],dataout_bnk3[3],dataout_bnk2[3],dataout_bnk1[3],dataout_bnk4[2],dataout_bnk3[2],dataout_bnk2[2],dataout_bnk1[2],dataout_bnk4[1],dataout_bnk3[1],dataout_bnk2[1],dataout_bnk1[1],dataout_bnk4[0],dataout_bnk3[0],dataout_bnk2[0],dataout_bnk1[0]}:{dataout_bnk4[15:0],dataout_bnk3[15:0],dataout_bnk2[15:0],dataout_bnk1[15:0] }) :
                 64'hxxxx_xxxx_xxxx_xxxx;			 
 
FIFOCTRL18KV1 # (
	.PEEK_MODE	(peek),
	.FIFO_EN	(1'b1),
	.R_WIDTH	(read_sel),
	.W_WIDTH	(write_sel),
	.DEPTH_EXT_MODE	({ext_18k, depth_extension}),
    .USR_PF     (prog_full),
	.USR_PE		(prog_empty)    
    )
u0_fifo_ctrl (
	.rst_n		(reset),
	.rd_req_n	(readen),
	.wr_req_n	(writeen),
	.clka		(readclk),
	.clkb		(writeclk),
	.write_drop	(writedrop),
	.write_save	(writesave),

	.full		(full),
	.empty		(empty),
	.prog_full	(almostfull),
	.prog_empty	(almostempty),
	.wptr		(wptr[13:0]),
	.rptr		(rptr[13:0]),
	.wr_mem_n	(wr_mem_n),
	.rd_mem_n	(rd_mem_n),
	.overflow	(overflow),
	.underflow	(underflow),
    .wrdp_rd_flag(writedropflag),
	.peek_en	(peek_en),
    .peek_rd_en (peek_rd_en)    
);

BRAM18KV1 # (
    .DEPTH_EXT_MODE23       (depth_extension),
    .DEPTH_EXT_MODE01       (depth_extension),
    .ECC_DEC_EN             (eccreaden),
    .ECC_ENC_EN             (eccwriteen),
    
    .EMB5K_4_MODEA_SEL      (read_sel),
    .EMB5K_4_MODEB_SEL      (write_sel),
    .EMB5K_4_PORTA_BYPASS   (1'b0),
    .EMB5K_4_PORTA_CE       (1'b1),
    .EMB5K_4_PORTA_REG_OUT  (outreg),
    .EMB5K_4_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_4_PORTA_CKINV    (readclk_inv),
    .EMB5K_4_PORTB_BYPASS   (1'b0),
    .EMB5K_4_PORTB_CE       (1'b1),
    .EMB5K_4_PORTB_REG_OUT  (outreg),
    .EMB5K_4_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_4_PORTB_CKINV    (writeclk_inv),
    
    .EMB5K_3_MODEA_SEL      (read_sel),
    .EMB5K_3_MODEB_SEL      (write_sel),
    .EMB5K_3_PORTA_BYPASS   (1'b0),
    .EMB5K_3_PORTA_CE       (1'b1),
    .EMB5K_3_PORTA_REG_OUT  (outreg),
    .EMB5K_3_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_3_PORTA_CKINV    (readclk_inv),
    .EMB5K_3_PORTB_BYPASS   (1'b0),
    .EMB5K_3_PORTB_CE       (1'b1),
    .EMB5K_3_PORTB_REG_OUT  (outreg),
    .EMB5K_3_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_3_PORTB_CKINV    (writeclk_inv),
    
    .EMB5K_2_MODEA_SEL      (read_sel),
    .EMB5K_2_MODEB_SEL      (write_sel),
    .EMB5K_2_PORTA_BYPASS   (1'b0),
    .EMB5K_2_PORTA_CE       (1'b1),
    .EMB5K_2_PORTA_REG_OUT  (outreg),
    .EMB5K_2_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_2_PORTA_CKINV    (readclk_inv),
    .EMB5K_2_PORTB_BYPASS   (1'b0),
    .EMB5K_2_PORTB_CE       (1'b1),
    .EMB5K_2_PORTB_REG_OUT  (outreg),
    .EMB5K_2_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_2_PORTB_CKINV    (writeclk_inv),
    
    .EMB5K_1_MODEA_SEL      (read_sel),
    .EMB5K_1_MODEB_SEL      (write_sel),
    .EMB5K_1_PORTA_BYPASS   (1'b0),
    .EMB5K_1_PORTA_CE       (1'b1),
    .EMB5K_1_PORTA_REG_OUT  (outreg),
    .EMB5K_1_PORTA_WR_MODE  (2'b01),    //write_first
    .EMB5K_1_PORTA_CKINV    (readclk_inv),
    .EMB5K_1_PORTB_BYPASS   (1'b0),
    .EMB5K_1_PORTB_CE       (1'b1),
    .EMB5K_1_PORTB_REG_OUT  (outreg),
    .EMB5K_1_PORTB_WR_MODE  (2'b01),    //write_first
    .EMB5K_1_PORTB_CKINV    (writeclk_inv),
    
    .EXT_18K                (ext_18k),
    .FIFO_EN                (1'b1),
    .PEEK_MODE              (peek),
    .PORTA_PROG             (8'b11110000),
    .PORTB_PROG             (8'b00001111),
    .WIDTH_EXT_MODE23       (width_extension),
    .WIDTH_EXT_MODE01       (width_extension)
    )
u0_emb18k_core (    
    .a_addr_ext             ({2'b11}),
    .b_addr_ext             ({2'b11}),
    
    .c1r4_aa                (),
    .c1r4_ab                (),
    .c1r4_cea               (),
    .c1r4_ceb               (),
    .c1r4_clka              (readclk),
    .c1r4_clkb              (writeclk),
    .c1r4_da                (),
    .c1r4_db                (datain_bnk4),
    .c1r4_rstna             (1'b1),
    .c1r4_rstnb             (1'b1),
    .c1r4_wea               (),
    .c1r4_web               (),
    .c1r4_user_ena          (regce),
    .c1r4_user_enb          (regce),
    
    .c1r3_aa                (),
    .c1r3_ab                (),
    .c1r3_cea               (),
    .c1r3_ceb               (),
    .c1r3_clka              (readclk),
    .c1r3_clkb              (writeclk),
    .c1r3_da                (),
    .c1r3_db                (datain_bnk3),
    .c1r3_rstna             (1'b1),
    .c1r3_rstnb             (1'b1),
    .c1r3_wea               (),
    .c1r3_web               (),
    .c1r3_user_ena          (regce),
    .c1r3_user_enb          (regce),
    
    .c1r2_aa                (),
    .c1r2_ab                (),
    .c1r2_cea               (),
    .c1r2_ceb               (),
    .c1r2_clka              (readclk),
    .c1r2_clkb              (writeclk),
    .c1r2_da                (),
    .c1r2_db                (datain_bnk2),
    .c1r2_rstna             (1'b1),
    .c1r2_rstnb             (1'b1),
    .c1r2_wea               (),
    .c1r2_web               (),
    .c1r2_user_ena          (regce),
    .c1r2_user_enb          (regce),    
    
    .c1r1_aa                (),
    .c1r1_ab                (),
    .c1r1_cea               (),
    .c1r1_ceb               (),
    .c1r1_clka              (readclk),
    .c1r1_clkb              (writeclk),
    .c1r1_da                (),
    .c1r1_db                (datain_bnk1),
    .c1r1_rstna             (reset),
    .c1r1_rstnb             (1'b1),
    .c1r1_wea               (),
    .c1r1_web               (),
    .c1r1_user_ena          (regce),
    .c1r1_user_enb          (regce),
    
    .rd_mem_n               (rd_mem_n),
    .rptr                   (rptr[13:0]),
    .wptr                   (wptr[13:0]),
    .wr_mem_n               (wr_mem_n),
    .peek_en                (peek_en),
    .peek_rd_en             (peek_rd_en),
        
    .c1r4_q                 (dataout_bnk4),
    .c1r3_q                 (dataout_bnk3),
    .c1r2_q                 (dataout_bnk2),
    .c1r1_q                 (dataout_bnk1),
    .eccindberr		        (eccindberr),
    .eccinsberr		        (eccinsberr),
    .eccoutdberr	        (eccoutdberr),
    .eccoutsberr	        (eccoutsberr),
    .err_addr		        (eccreadaddr) 
);     
    
endmodule // FIFO18K

// end of FIFO18K 

module SIO (
    f_id,
    clk_en,
    fclk,
    od,
    oen,
    rstn,
    setn,
    PAD
);

input            clk_en;
input            fclk;
input    [1:0]    od;
input            oen;
input            rstn;
input            setn;

output    [1:0]    f_id;

inout            PAD;

//Analog IO parameters
parameter   KEEP      = 2'b0;
parameter   NDR       = 4'b0;
parameter   NS_LV     = 2'b0;
parameter   PDR       = 4'b0;
parameter   RX_DIG_EN = 1'b0;
parameter   VPCI_EN   = 1'b0;

//Logic IO/IOC parameters
parameter   OEN_SEL      = 2'b0;    //2'b00 :  1'b1
                                    //2'b01 :  1'b0
                                    //2'b10 :  f_oen
                                    //2'b11 : ~f_oen
parameter   OUT_SEL      = 2'b0;    //2'b00 :  1'b1
                                    //2'b01 :  1'b0
                                    //2'b10 :  f_od
                                    //2'b11 : ~f_od

parameter   CLK_INV      = 1'b0;    //1'b1 : ~fclk
                                    //1'b0 : fclk
parameter   FCLK_GATE_EN = 1'b0;    //1'b0 : no clock gating
                                    //1'b1 : clock gating use clk_en
parameter   SETN_INV     = 1'b0;    //1'b1 : setn inverted
                                    //1'b0 : setn not inverted
parameter   SETN_SYNC    = 1'b0;    //1'b1 : setn sync
                                    //1'b0 : setn async
parameter   RSTN_INV     = 1'b0;    //1'b1 : rstn inverted
                                    //1'b0 : rstn not inverted
parameter   RSTN_SYNC    = 1'b0;    //1'b1 : rstn sync
                                    //1'b0 : rstn async
parameter   OEN_SETN_EN  = 1'b0;    //1'b1 : oen setn enabled
                                    //1'b0 : oen setn disabled
parameter   OD_SETN_EN   = 1'b0;    //1'b1 : od setn enabled
                                    //1'b0 : od setn disabled
parameter   ID_SETN_EN   = 1'b0;    //1'b1 : id setn enabled
                                    //1'b0 : id setn disabled
parameter   OEN_RSTN_EN  = 1'b0;    //1'b1 : oen rstn enabled
                                    //1'b0 : oen rstn disabled
parameter   OD_RSTN_EN   = 1'b0;    //1'b1 : od rstn enabled
                                    //1'b0 : od rstn disabled
parameter   ID_RSTN_EN   = 1'b0;    //1'b1 : id rstn enabled
                                    //1'b0 : id rstn disabled
parameter   FOEN_SEL    = 1'b0;     //1'b1 : registered
                                    //1'b0 : bypassed
parameter   FOUT_SEL    = 1'b0;     //1'b1 : registered
                                    //1'b0 : bypassed
parameter   FIN_SEL     = 1'b0;     //1'b1 : registered
                                    //1'b0 : bypassed
parameter   DDR_EN       = 1'b0;    //DDR enable
parameter   DDR_REG_EN   = 1'b0;    //SDR fast output: DDR_REG = 1'b0 && FOUT_SEL = 1'b1
                                    //DDR with 1 pipeline: DDR_REG = 1'b1 && FOUT_SEL = 1'b1
parameter   DDR_PREG_EN  = 1'b0;    //SDR fast input: DDR_PREG = 1'b0 && FIN_SEL = 1'b1
                                    //DDR with 1 pipeline: DDR_PREG = 1'b1 && FOUT_SEL = 1'b1
parameter   DDR_NREG_EN  = 1'b0;

parameter   is_clk_io = "false";
parameter   optional_function = ""; //"spi_sclk", "spi_sdi", "spi_cson", "spi_sdo", "spi_wpn", "spi_holdn"

wire        f_od;
wire        f_oen;
wire        id;

BASIC_IO basic_io_inst0 (
    .f_od    (f_od),
    .f_oen    (f_oen),

    .id    (id),
    .PAD    (PAD)
);
defparam basic_io_inst0.CFG_KEEP      = KEEP;
defparam basic_io_inst0.CFG_NDR       = NDR;
defparam basic_io_inst0.CFG_NS_LV     = NS_LV;
defparam basic_io_inst0.CFG_PDR       = PDR;
defparam basic_io_inst0.CFG_RX_DIG_EN = RX_DIG_EN;
defparam basic_io_inst0.VPCI_EN       = VPCI_EN;

defparam basic_io_inst0.CFG_OEN_SEL   = OEN_SEL;
defparam basic_io_inst0.CFG_OUT_SEL   = OUT_SEL;

IOC_CMOS ioc_cmos_inst0 (
    .clk_en    (clk_en),
    .fclk    (fclk),
    .id    (id),
    .od    (od[1:0]),
    .oen    (oen),
    .rstn    (rstn),
    .setn    (setn),

    .f_id    (f_id[1:0]),
    .f_od    (f_od),
    .f_oen    (f_oen)
);
defparam ioc_cmos_inst0.CFG_CLK_INV      = CLK_INV;
defparam ioc_cmos_inst0.CFG_FCLK_GATE_EN = FCLK_GATE_EN;
defparam ioc_cmos_inst0.CFG_SETN_INV     = SETN_INV;
defparam ioc_cmos_inst0.CFG_SETN_SYNC    = SETN_SYNC;
defparam ioc_cmos_inst0.CFG_OEN_SETN_EN  = OEN_SETN_EN;
defparam ioc_cmos_inst0.CFG_OD_SETN_EN   = OD_SETN_EN;
defparam ioc_cmos_inst0.CFG_ID_SETN_EN   = ID_SETN_EN;
defparam ioc_cmos_inst0.CFG_RSTN_INV     = RSTN_INV;
defparam ioc_cmos_inst0.CFG_RSTN_SYNC    = RSTN_SYNC;
defparam ioc_cmos_inst0.CFG_OEN_RSTN_EN  = OEN_RSTN_EN;
defparam ioc_cmos_inst0.CFG_OD_RSTN_EN   = OD_RSTN_EN;
defparam ioc_cmos_inst0.CFG_ID_RSTN_EN   = ID_RSTN_EN;
defparam ioc_cmos_inst0.CFG_FOEN_SELN    = !FOEN_SEL;
defparam ioc_cmos_inst0.CFG_FOUT_SELN    = !FOUT_SEL;
defparam ioc_cmos_inst0.CFG_FIN_SELN     = !FIN_SEL;
defparam ioc_cmos_inst0.CFG_DDR          = DDR_EN;
defparam ioc_cmos_inst0.CFG_DDR_REG      = DDR_REG_EN;
defparam ioc_cmos_inst0.CFG_DDR_PREG     = DDR_PREG_EN;
defparam ioc_cmos_inst0.CFG_DDR_NREG     = DDR_NREG_EN;

endmodule

//For EMB_Wizard Begin
module CS_REG_PRIM(Q, D, CLK, RST, SET, CE);
 
   output Q;
   input  D, CLK, RST, SET, CE;
 
   wire                 INIT = 1'bX;
   reg                  QX_REG;
 
   initial begin
      QX_REG = INIT;
   end
 
 
   wire SET_PRI = SET && !RST;       // Force priority
 
   always @(posedge CLK) begin
      if (CE) begin
              if (RST) QX_REG <= 1'b0;
                  else if (SET) QX_REG <= 1'b1;
                  else QX_REG <= D;
          end
   end
 
   assign Q = QX_REG;
 
endmodule

module CS_GND_PRIM(OUT);

   output        OUT;
   parameter        PLACE_LOCATION = "NONE";
   parameter        PCK_LOCATION = "NONE";


   assign         OUT = 1'b0;

endmodule

module CS_VCC_PRIM(OUT);

   output        OUT;
   parameter        PLACE_LOCATION = "NONE";
   parameter        PCK_LOCATION = "NONE";

   assign         OUT = 1'b1;
   
endmodule

module CS_REG_E_PRIM(Q, D, CLK, CE);

   output Q;
   input  D, CLK, CE;

wire gnd_inst;

CS_GND_PRIM gnd (
    .OUT(gnd_inst)
);
   
CS_REG_PRIM reg_r (
    .CLK(CLK ), 
    .D(D ), 
    .Q(Q ), 
    .RST(gnd_inst ),
    .SET(gnd_inst ),
    .CE(CE )
);   
endmodule

module CS_REG_CLK_PRIM(Q, D, CLK);

   output Q;
   input  D, CLK;

wire vcc_inst;
wire gnd_inst;

CS_VCC_PRIM vcc (
    .OUT(vcc_inst)
);

CS_GND_PRIM gnd (
    .OUT(gnd_inst)
);
   
CS_REG_PRIM reg_r (
    .CLK(CLK ), 
    .D(D ), 
    .Q(Q ), 
    .RST(gnd_inst ),
    .SET(gnd_inst ),
    .CE(vcc_inst )
);   
endmodule

module mx2a(Y, D0, D1, S);
        input D0;
        input D1;
        input S;
        output Y;

    assign Y = (!S&D0)|(S&D1);
endmodule

module CS_BUF_PRIM (A, Y);
        input A;
        output Y;

    assign Y = A;
endmodule

module CS_INV_PRIM (OUT, IN);

   output  OUT;    
   input   IN;    
   parameter        PLACE_LOCATION = "NONE";
   parameter        PCK_LOCATION = "NONE";
   
   assign    OUT = !IN;
 
endmodule

module AND2 (O, I0, I1);
        input I0;
        input I1;
        output O;

    assign O = I1&I0;
endmodule

//For EMB_Wizard End

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////


module ADC (
    fp_adc_int_o,
    fp_adc_pbus_gnt,
    fp_adc_pbus_rdata,
    fp_adc_pbus_addr,
    fp_adc_pbus_req,
    fp_adc_pbus_wdata,
    fp_adc_pbus_write,
    fp_clk_adc,
    fp_rst_adc_n,
    ana_ADC_ADION,
    ana_ADC_ADIOP,
    ana_ADC_VINN,
    ana_ADC_VINP,
    ana_ADC_VIPN,
    ana_ADC_VIPP,
    ana_ADC_VREFN,
    ana_ADC_VREFP
);

//Connection with FP
output             fp_adc_int_o;
output             fp_adc_pbus_gnt;
output    [31:0]   fp_adc_pbus_rdata;
input    [7:0]     fp_adc_pbus_addr;
input              fp_adc_pbus_req;
input    [31:0]    fp_adc_pbus_wdata;
input              fp_adc_pbus_write;
input              fp_clk_adc;
input              fp_rst_adc_n;

//PADS
input    [11:0]    ana_ADC_ADION;              //share digital input pairs
input    [11:0]    ana_ADC_ADIOP;              //share digital input pairs
input              ana_ADC_VINN;               //analog input pairs
input              ana_ADC_VINP;               //analog input pairs
input              ana_ADC_VIPN;               //analog input pairs
input              ana_ADC_VIPP;               //analog input pairs
inout              ana_ADC_VREFN;              //vrefn
inout              ana_ADC_VREFP;              //vrefp

parameter   adc_amux_sel   = 2'b00;   //[5:4]
parameter   adc_bg_pd      = 1'b1;    //[3]
parameter   adc_cf_fp_sel  = 1'b0;    //[0]
parameter   adc_clk_gate   = 1'b0;    //[2]
parameter   adc_clk_inv    = 1'b1;    //[1]

endmodule

// 1-bit full adder
//------------------------------------
module ADD_1BIT (
	s,
	co,
	p,
	pb,
	
	ci,
	b,
	a
);

output     s;
output     co;
output     p;
output     pb;

input      ci;
input      b;
input      a;

`ifndef CS_SW_SKEL
    assign p  = a ^ b;
    assign pb = ~p;
    assign co = p ? ci : a ;
    assign s  = ci ^ p;

specify

   (ci => co)   = (0,0);
   (a  => co)   = (0,0);
   (b  => co)   = (0,0);

   (ci => s)    = (0,0);
   (a  => s)    = (0,0);
   (b  => s)    = (0,0);

   (a  => p)    = (0,0);
   (b  => p)    = (0,0);

   (a  => pb)   = (0,0);
   (b  => pb)   = (0,0);
            
endspecify
    
`endif



endmodule

module AND4 (
	o,
	
	a,
	b,
	c,
	d
	);

output	o;

input a;
input b;
input c;
input d;

`ifndef CS_SW_SKEL
    assign    o = (a & b) & (c & d);
    
    specify

    ( a => o ) = (0,0);
    ( b => o ) = (0,0);
    ( c => o ) = (0,0);
    ( d => o ) = (0,0);

    endspecify
`endif

endmodule
module BASIC_IO(
	 id
	,f_od
	,f_oen
	,PAD
`ifdef FM_HACK
	,CFG_KEEP
	,CFG_NDR
	,CFG_NS_LV
	,CFG_OEN_SEL
	,CFG_OUT_SEL
	,CFG_PDR
	,CFG_RX_DIG_EN
	,VPCI_EN
`endif
);

output		id;
input		f_od;
input		f_oen;
inout		PAD;
`ifdef FM_HACK
input	[1:0]	CFG_KEEP;
input	[3:0]	CFG_NDR;
input	[1:0]	CFG_NS_LV;
input	[1:0]	CFG_OEN_SEL;
input	[1:0]	CFG_OUT_SEL;
input	[3:0]	CFG_PDR;
input		CFG_RX_DIG_EN;
input		VPCI_EN;
`else
parameter 	CFG_KEEP         = 2'b0;
parameter 	CFG_NDR          = 4'b0;
parameter 	CFG_NS_LV        = 2'b0;
parameter 	CFG_OEN_SEL      = 2'b0;
parameter 	CFG_OUT_SEL      = 2'b0;
parameter 	CFG_PDR          = 4'b0;
parameter 	CFG_RX_DIG_EN    = 1'b0;
parameter 	VPCI_EN          = 1'b0;
`endif

io_data data_path (
	.f_oen		(f_oen),
	.f_od		(f_od),
	.rxd		(RXD),
	.CFG_OEN_SEL	(CFG_OEN_SEL[1:0]),
	.CFG_OUT_SEL	(CFG_OUT_SEL[1:0]),

	.id		(id),
	.ted		(TED),
	.txd		(TXD) 
);

CSGPIO ana_IO (
	.TXD		(TXD),
	.TED		(TED),
	.NS_LV		(CFG_NS_LV[1:0]),
	.PDR		(CFG_PDR[3:0]),
	.NDR		(CFG_NDR[3:0]),
	.KEEP		(CFG_KEEP[1:0]),
	.RX_DIG_EN	(CFG_RX_DIG_EN),
	.VPCI_EN	(VPCI_EN),

	.RXD		(RXD),
	.PAD		(PAD)
);

endmodule


// VPERL: GENERATED_BEG

module BRAM18KV1 (
	c1r4_q,
	c1r3_q,
	c1r2_q,
	c1r1_q,
	eccoutdberr,
	eccoutsberr,
	err_addr,
	a_addr_ext,
	b_addr_ext,
	c1r4_aa,
	c1r4_ab,
	c1r4_cea,
	c1r4_ceb,
	c1r4_clka,
	c1r4_clkb,
	c1r4_da,
	c1r4_db,
	c1r4_rstna,
	c1r4_rstnb,
	c1r4_user_ena,
	c1r4_user_enb,
	c1r4_wea,
	c1r4_web,
	c1r3_aa,
	c1r3_ab,
	c1r3_cea,
	c1r3_ceb,
	c1r3_clka,
	c1r3_clkb,
	c1r3_da,
	c1r3_db,
	c1r3_rstna,
	c1r3_rstnb,
	c1r3_user_ena,
	c1r3_user_enb,
	c1r3_wea,
	c1r3_web,
	c1r2_aa,
	c1r2_ab,
	c1r2_cea,
	c1r2_ceb,
	c1r2_clka,
	c1r2_clkb,
	c1r2_da,
	c1r2_db,
	c1r2_rstna,
	c1r2_rstnb,
	c1r2_user_ena,
	c1r2_user_enb,
	c1r2_wea,
	c1r2_web,
	c1r1_aa,
	c1r1_ab,
	c1r1_cea,
	c1r1_ceb,
	c1r1_clka,
	c1r1_clkb,
	c1r1_da,
	c1r1_db,
	c1r1_rstna,
	c1r1_rstnb,
	c1r1_user_ena,
	c1r1_user_enb,
	c1r1_wea,
	c1r1_web,
	eccindberr,
	eccinsberr,
	peek_en,
	peek_rd_en,
	rd_mem_n,
	rptr,
	wptr,
	wr_mem_n 
`ifdef FM_HACK
    ,DEC_REG_EN
    ,DEPTH_EXT_MODE23
    ,DEPTH_EXT_MODE01
    ,ECC_DEC_EN
    ,ECC_ENC_EN
    ,EMB5K_4_MODEA_SEL
    ,EMB5K_4_MODEB_SEL
    ,EMB5K_4_PORTA_BYPASS
    ,EMB5K_4_PORTA_CE
    ,EMB5K_4_PORTA_CKINV
    ,EMB5K_4_PORTA_REG_OUT
    ,EMB5K_4_PORTA_WR_MODE
    ,EMB5K_4_PORTB_BYPASS
    ,EMB5K_4_PORTB_CE
    ,EMB5K_4_PORTB_CKINV
    ,EMB5K_4_PORTB_REG_OUT
    ,EMB5K_4_PORTB_WR_MODE
    ,EMB5K_3_MODEA_SEL
    ,EMB5K_3_MODEB_SEL
    ,EMB5K_3_PORTA_BYPASS
    ,EMB5K_3_PORTA_CE
    ,EMB5K_3_PORTA_CKINV
    ,EMB5K_3_PORTA_REG_OUT
    ,EMB5K_3_PORTA_WR_MODE
    ,EMB5K_3_PORTB_BYPASS
    ,EMB5K_3_PORTB_CE
    ,EMB5K_3_PORTB_CKINV
    ,EMB5K_3_PORTB_REG_OUT
    ,EMB5K_3_PORTB_WR_MODE
    ,EMB5K_2_MODEA_SEL
    ,EMB5K_2_MODEB_SEL
    ,EMB5K_2_PORTA_BYPASS
    ,EMB5K_2_PORTA_CE
    ,EMB5K_2_PORTA_CKINV
    ,EMB5K_2_PORTA_REG_OUT
    ,EMB5K_2_PORTA_WR_MODE
    ,EMB5K_2_PORTB_BYPASS
    ,EMB5K_2_PORTB_CE
    ,EMB5K_2_PORTB_CKINV
    ,EMB5K_2_PORTB_REG_OUT
    ,EMB5K_2_PORTB_WR_MODE
    ,EMB5K_1_MODEA_SEL
    ,EMB5K_1_MODEB_SEL
    ,EMB5K_1_PORTA_BYPASS
    ,EMB5K_1_PORTA_CE
    ,EMB5K_1_PORTA_CKINV
    ,EMB5K_1_PORTA_REG_OUT
    ,EMB5K_1_PORTA_WR_MODE
    ,EMB5K_1_PORTB_BYPASS
    ,EMB5K_1_PORTB_CE
    ,EMB5K_1_PORTB_CKINV
    ,EMB5K_1_PORTB_REG_OUT
    ,EMB5K_1_PORTB_WR_MODE
    ,EXT_18K
    ,FIFO_EN
    ,PEEK_MODE
    ,PORTA_PROG
    ,PORTB_PROG
    ,WIDTH_EXT_MODE23
    ,WIDTH_EXT_MODE01
`endif
);

output	[17:0]	c1r4_q;
output	[17:0]	c1r3_q;
output	[17:0]	c1r2_q;
output	[17:0]	c1r1_q;
output		eccoutdberr;
output		eccoutsberr;
output	[7:0]	err_addr;
input	[1:0]	a_addr_ext;
input	[1:0]	b_addr_ext;
input	[11:0]	c1r4_aa;
input	[11:0]	c1r4_ab;
input		c1r4_cea;
input		c1r4_ceb;
input		c1r4_clka;
input		c1r4_clkb;
input	[17:0]	c1r4_da;
input	[17:0]	c1r4_db;
input		c1r4_rstna;
input		c1r4_rstnb;
input		c1r4_user_ena;
input		c1r4_user_enb;
input		c1r4_wea;
input		c1r4_web;
input	[11:0]	c1r3_aa;
input	[11:0]	c1r3_ab;
input		c1r3_cea;
input		c1r3_ceb;
input		c1r3_clka;
input		c1r3_clkb;
input	[17:0]	c1r3_da;
input	[17:0]	c1r3_db;
input		c1r3_rstna;
input		c1r3_rstnb;
input		c1r3_user_ena;
input		c1r3_user_enb;
input		c1r3_wea;
input		c1r3_web;
input	[11:0]	c1r2_aa;
input	[11:0]	c1r2_ab;
input		c1r2_cea;
input		c1r2_ceb;
input		c1r2_clka;
input		c1r2_clkb;
input	[17:0]	c1r2_da;
input	[17:0]	c1r2_db;
input		c1r2_rstna;
input		c1r2_rstnb;
input		c1r2_user_ena;
input		c1r2_user_enb;
input		c1r2_wea;
input		c1r2_web;
input	[11:0]	c1r1_aa;
input	[11:0]	c1r1_ab;
input		c1r1_cea;
input		c1r1_ceb;
input		c1r1_clka;
input		c1r1_clkb;
input	[17:0]	c1r1_da;
input	[17:0]	c1r1_db;
input		c1r1_rstna;
input		c1r1_rstnb;
input		c1r1_user_ena;
input		c1r1_user_enb;
input		c1r1_wea;
input		c1r1_web;
input		eccindberr;
input		eccinsberr;
input		peek_en;
input		peek_rd_en;
input		rd_mem_n;
input	[13:0]	rptr;
input	[13:0]	wptr;
input		wr_mem_n;

`ifdef FM_HACK
input         DEC_REG_EN;
input         DEPTH_EXT_MODE23;
input         DEPTH_EXT_MODE01;
input         ECC_DEC_EN;
input         ECC_ENC_EN;
input  [3:0]  EMB5K_4_MODEA_SEL;
input  [3:0]  EMB5K_4_MODEB_SEL;
input         EMB5K_4_PORTA_BYPASS;
input         EMB5K_4_PORTA_CE;
input         EMB5K_4_PORTA_CKINV;
input         EMB5K_4_PORTA_REG_OUT;
input  [1:0]  EMB5K_4_PORTA_WR_MODE;
input         EMB5K_4_PORTB_BYPASS;
input         EMB5K_4_PORTB_CE;
input         EMB5K_4_PORTB_CKINV;
input         EMB5K_4_PORTB_REG_OUT;
input  [1:0]  EMB5K_4_PORTB_WR_MODE;
input  [3:0]  EMB5K_3_MODEA_SEL;
input  [3:0]  EMB5K_3_MODEB_SEL;
input         EMB5K_3_PORTA_BYPASS;
input         EMB5K_3_PORTA_CE;
input         EMB5K_3_PORTA_CKINV;
input         EMB5K_3_PORTA_REG_OUT;
input  [1:0]  EMB5K_3_PORTA_WR_MODE;
input         EMB5K_3_PORTB_BYPASS;
input         EMB5K_3_PORTB_CE;
input         EMB5K_3_PORTB_CKINV;
input         EMB5K_3_PORTB_REG_OUT;
input  [1:0]  EMB5K_3_PORTB_WR_MODE;
input  [3:0]  EMB5K_2_MODEA_SEL;
input  [3:0]  EMB5K_2_MODEB_SEL;
input         EMB5K_2_PORTA_BYPASS;
input         EMB5K_2_PORTA_CE;
input         EMB5K_2_PORTA_CKINV;
input         EMB5K_2_PORTA_REG_OUT;
input  [1:0]  EMB5K_2_PORTA_WR_MODE;
input         EMB5K_2_PORTB_BYPASS;
input         EMB5K_2_PORTB_CE;
input         EMB5K_2_PORTB_CKINV;
input         EMB5K_2_PORTB_REG_OUT;
input  [1:0]  EMB5K_2_PORTB_WR_MODE;
input  [3:0]  EMB5K_1_MODEA_SEL;
input  [3:0]  EMB5K_1_MODEB_SEL;
input         EMB5K_1_PORTA_BYPASS;
input         EMB5K_1_PORTA_CE;
input         EMB5K_1_PORTA_CKINV;
input         EMB5K_1_PORTA_REG_OUT;
input  [1:0]  EMB5K_1_PORTA_WR_MODE;
input         EMB5K_1_PORTB_BYPASS;
input         EMB5K_1_PORTB_CE;
input         EMB5K_1_PORTB_CKINV;
input         EMB5K_1_PORTB_REG_OUT;
input  [1:0]  EMB5K_1_PORTB_WR_MODE;
input         EXT_18K;
input         FIFO_EN;
input         PEEK_MODE;
input  [7:0]  PORTA_PROG;
input  [7:0]  PORTB_PROG;
input         WIDTH_EXT_MODE23;
input         WIDTH_EXT_MODE01;
`else
parameter                DEC_REG_EN                               = 1'b0;
parameter                DEPTH_EXT_MODE23                         = 1'b0;
parameter                DEPTH_EXT_MODE01                         = 1'b0;
parameter                ECC_DEC_EN                               = 1'b0;
parameter                ECC_ENC_EN                               = 1'b0;
parameter                EMB5K_4_MODEA_SEL                        = 4'b0;
parameter                EMB5K_4_MODEB_SEL                        = 4'b0;
parameter                EMB5K_4_PORTA_BYPASS                     = 1'b0;
parameter                EMB5K_4_PORTA_CE                         = 1'b0;
parameter                EMB5K_4_PORTA_CKINV                      = 1'b0;
parameter                EMB5K_4_PORTA_REG_OUT                    = 1'b0;
parameter                EMB5K_4_PORTA_WR_MODE                    = 2'b0;
parameter                EMB5K_4_PORTB_BYPASS                     = 1'b0;
parameter                EMB5K_4_PORTB_CE                         = 1'b0;
parameter                EMB5K_4_PORTB_CKINV                      = 1'b0;
parameter                EMB5K_4_PORTB_REG_OUT                    = 1'b0;
parameter                EMB5K_4_PORTB_WR_MODE                    = 2'b0;
parameter                EMB5K_3_MODEA_SEL                        = 4'b0;
parameter                EMB5K_3_MODEB_SEL                        = 4'b0;
parameter                EMB5K_3_PORTA_BYPASS                     = 1'b0;
parameter                EMB5K_3_PORTA_CE                         = 1'b0;
parameter                EMB5K_3_PORTA_CKINV                      = 1'b0;
parameter                EMB5K_3_PORTA_REG_OUT                    = 1'b0;
parameter                EMB5K_3_PORTA_WR_MODE                    = 2'b0;
parameter                EMB5K_3_PORTB_BYPASS                     = 1'b0;
parameter                EMB5K_3_PORTB_CE                         = 1'b0;
parameter                EMB5K_3_PORTB_CKINV                      = 1'b0;
parameter                EMB5K_3_PORTB_REG_OUT                    = 1'b0;
parameter                EMB5K_3_PORTB_WR_MODE                    = 2'b0;
parameter                EMB5K_2_MODEA_SEL                        = 4'b0;
parameter                EMB5K_2_MODEB_SEL                        = 4'b0;
parameter                EMB5K_2_PORTA_BYPASS                     = 1'b0;
parameter                EMB5K_2_PORTA_CE                         = 1'b0;
parameter                EMB5K_2_PORTA_CKINV                      = 1'b0;
parameter                EMB5K_2_PORTA_REG_OUT                    = 1'b0;
parameter                EMB5K_2_PORTA_WR_MODE                    = 2'b0;
parameter                EMB5K_2_PORTB_BYPASS                     = 1'b0;
parameter                EMB5K_2_PORTB_CE                         = 1'b0;
parameter                EMB5K_2_PORTB_CKINV                      = 1'b0;
parameter                EMB5K_2_PORTB_REG_OUT                    = 1'b0;
parameter                EMB5K_2_PORTB_WR_MODE                    = 2'b0;
parameter                EMB5K_1_MODEA_SEL                        = 4'b0;
parameter                EMB5K_1_MODEB_SEL                        = 4'b0;
parameter                EMB5K_1_PORTA_BYPASS                     = 1'b0;
parameter                EMB5K_1_PORTA_CE                         = 1'b0;
parameter                EMB5K_1_PORTA_CKINV                      = 1'b0;
parameter                EMB5K_1_PORTA_REG_OUT                    = 1'b0;
parameter                EMB5K_1_PORTA_WR_MODE                    = 2'b0;
parameter                EMB5K_1_PORTB_BYPASS                     = 1'b0;
parameter                EMB5K_1_PORTB_CE                         = 1'b0;
parameter                EMB5K_1_PORTB_CKINV                      = 1'b0;
parameter                EMB5K_1_PORTB_REG_OUT                    = 1'b0;
parameter                EMB5K_1_PORTB_WR_MODE                    = 2'b0;
parameter                EXT_18K                                  = 1'b0;
parameter                FIFO_EN                                  = 1'b0;
parameter                PEEK_MODE                                = 1'b0;
parameter                PORTA_PROG                               = 8'b0;
parameter                PORTB_PROG                               = 8'b0;
parameter                WIDTH_EXT_MODE23                         = 1'b0;
parameter                WIDTH_EXT_MODE01                         = 1'b0;
`endif

`ifndef FM_HACK
    reg gbl_clear_b=1;
    wire GSR;
    glbsr inst( .GSR( GSR )) ;

    initial begin
        gbl_clear_b = 1'b0;
        @(posedge GSR);
        gbl_clear_b = 1'b1;
    end

    parameter init_00_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

    parameter init_00_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

    parameter init_00_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    
    parameter init_00_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_01_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_02_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_03_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_04_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_05_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_06_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_07_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_08_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_09_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0a_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0b_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0c_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0d_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0e_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter init_0f_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_00_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter initp_01_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

    initial begin
        force c1r1_rstna = 1'b0;
        force c1r1_rstnb = 1'b0;
        force c1r2_rstna = 1'b0;
        force c1r2_rstnb = 1'b0;
        force c1r3_rstna = 1'b0;
        force c1r3_rstnb = 1'b0;
        force c1r4_rstna = 1'b0;
        force c1r4_rstnb = 1'b0;
        @(posedge GSR);
        release c1r1_rstna;
        release c1r1_rstnb;
        release c1r2_rstna;
        release c1r2_rstnb;
        release c1r3_rstna;
        release c1r3_rstnb;
        release c1r4_rstna;
        release c1r4_rstnb;
    end

    integer i;
/*
    initial
    begin
    @(posedge GSR);
        for (i = 0; i < 16; i = i + 1)
        begin
            emb5k_core_1.emb5k_top.mem[i    ] <= {initp_00_1[i*2+1   -:2 ], init_00_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+16 ] <= {initp_00_1[i*2+33  -:2 ], init_01_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+32 ] <= {initp_00_1[i*2+65  -:2 ], init_02_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+48 ] <= {initp_00_1[i*2+97  -:2 ], init_03_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+64 ] <= {initp_00_1[i*2+129 -:2 ], init_04_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+80 ] <= {initp_00_1[i*2+161 -:2 ], init_05_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+96 ] <= {initp_00_1[i*2+193 -:2 ], init_06_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+112] <= {initp_00_1[i*2+225 -:2 ], init_07_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+128] <= {initp_01_1[i*2+1   -:2 ], init_08_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+144] <= {initp_01_1[i*2+33  -:2 ], init_09_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+160] <= {initp_01_1[i*2+65  -:2 ], init_0a_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+176] <= {initp_01_1[i*2+97  -:2 ], init_0b_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+192] <= {initp_01_1[i*2+129 -:2 ], init_0c_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+208] <= {initp_01_1[i*2+161 -:2 ], init_0d_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+224] <= {initp_01_1[i*2+193 -:2 ], init_0e_1[i*16+15 -:16 ]};
            emb5k_core_1.emb5k_top.mem[i+240] <= {initp_01_1[i*2+225 -:2 ], init_0f_1[i*16+15 -:16 ]};
        end
    end
    
    initial
    begin
    @(posedge GSR);
        for (i = 0; i < 16; i = i + 1)
        begin
            emb5k_core_2.emb5k_top.mem[i    ] <= {initp_00_2[i*2+1   -:2 ], init_00_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+16 ] <= {initp_00_2[i*2+33  -:2 ], init_01_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+32 ] <= {initp_00_2[i*2+65  -:2 ], init_02_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+48 ] <= {initp_00_2[i*2+97  -:2 ], init_03_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+64 ] <= {initp_00_2[i*2+129 -:2 ], init_04_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+80 ] <= {initp_00_2[i*2+161 -:2 ], init_05_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+96 ] <= {initp_00_2[i*2+193 -:2 ], init_06_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+112] <= {initp_00_2[i*2+225 -:2 ], init_07_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+128] <= {initp_01_2[i*2+1   -:2 ], init_08_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+144] <= {initp_01_2[i*2+33  -:2 ], init_09_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+160] <= {initp_01_2[i*2+65  -:2 ], init_0a_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+176] <= {initp_01_2[i*2+97  -:2 ], init_0b_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+192] <= {initp_01_2[i*2+129 -:2 ], init_0c_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+208] <= {initp_01_2[i*2+161 -:2 ], init_0d_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+224] <= {initp_01_2[i*2+193 -:2 ], init_0e_2[i*16+15 -:16 ]};
            emb5k_core_2.emb5k_top.mem[i+240] <= {initp_01_2[i*2+225 -:2 ], init_0f_2[i*16+15 -:16 ]};
        end
    end
    
    initial
    begin
    @(posedge GSR);
        for (i = 0; i < 16; i = i + 1)
        begin
            emb5k_core_3.emb5k_top.mem[i    ] <= {initp_00_3[i*2+1   -:2 ], init_00_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+16 ] <= {initp_00_3[i*2+33  -:2 ], init_01_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+32 ] <= {initp_00_3[i*2+65  -:2 ], init_02_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+48 ] <= {initp_00_3[i*2+97  -:2 ], init_03_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+64 ] <= {initp_00_3[i*2+129 -:2 ], init_04_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+80 ] <= {initp_00_3[i*2+161 -:2 ], init_05_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+96 ] <= {initp_00_3[i*2+193 -:2 ], init_06_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+112] <= {initp_00_3[i*2+225 -:2 ], init_07_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+128] <= {initp_01_3[i*2+1   -:2 ], init_08_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+144] <= {initp_01_3[i*2+33  -:2 ], init_09_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+160] <= {initp_01_3[i*2+65  -:2 ], init_0a_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+176] <= {initp_01_3[i*2+97  -:2 ], init_0b_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+192] <= {initp_01_3[i*2+129 -:2 ], init_0c_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+208] <= {initp_01_3[i*2+161 -:2 ], init_0d_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+224] <= {initp_01_3[i*2+193 -:2 ], init_0e_3[i*16+15 -:16 ]};
            emb5k_core_3.emb5k_top.mem[i+240] <= {initp_01_3[i*2+225 -:2 ], init_0f_3[i*16+15 -:16 ]};
        end
    end
    
    initial
    begin
    @(posedge GSR);
        for (i = 0; i < 16; i = i + 1)
        begin
            emb5k_core_4.emb5k_top.mem[i    ] <= {initp_00_4[i*2+1   -:2 ], init_00_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+16 ] <= {initp_00_4[i*2+33  -:2 ], init_01_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+32 ] <= {initp_00_4[i*2+65  -:2 ], init_02_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+48 ] <= {initp_00_4[i*2+97  -:2 ], init_03_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+64 ] <= {initp_00_4[i*2+129 -:2 ], init_04_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+80 ] <= {initp_00_4[i*2+161 -:2 ], init_05_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+96 ] <= {initp_00_4[i*2+193 -:2 ], init_06_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+112] <= {initp_00_4[i*2+225 -:2 ], init_07_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+128] <= {initp_01_4[i*2+1   -:2 ], init_08_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+144] <= {initp_01_4[i*2+33  -:2 ], init_09_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+160] <= {initp_01_4[i*2+65  -:2 ], init_0a_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+176] <= {initp_01_4[i*2+97  -:2 ], init_0b_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+192] <= {initp_01_4[i*2+129 -:2 ], init_0c_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+208] <= {initp_01_4[i*2+161 -:2 ], init_0d_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+224] <= {initp_01_4[i*2+193 -:2 ], init_0e_4[i*16+15 -:16 ]};
            emb5k_core_4.emb5k_top.mem[i+240] <= {initp_01_4[i*2+225 -:2 ], init_0f_4[i*16+15 -:16 ]};
        end
    end
*/
`else
    wire gbl_clear_b = 1;
`endif

wire	[11:0]	c1r4_aa_t;
wire	[11:0]	c1r4_ab_t;
wire		c1r4_cea_t;
wire		c1r4_ceb_t;
wire		c1r4_clka_inv;
wire		c1r4_clka_n;
wire		c1r4_clkb_inv;
wire		c1r4_clkb_n;
wire	[17:0]	c1r4_da_t;
wire	[17:0]	c1r4_db_ecc;
wire	[17:0]	c1r4_db_t;
wire	[17:0]	c1r4_q_t;
wire		c1r4_reg_ena;
wire		c1r4_reg_enb;
wire		c1r4_wea_t;
wire		c1r4_web_t;
wire	[11:0]	c1r3_aa_t;
wire	[11:0]	c1r3_ab_t;
wire		c1r3_cea_t;
wire		c1r3_ceb_t;
wire		c1r3_clka_inv;
wire		c1r3_clka_n;
wire		c1r3_clkb_inv;
wire		c1r3_clkb_n;
wire	[17:0]	c1r3_da_t;
wire	[17:0]	c1r3_db_ecc;
wire	[17:0]	c1r3_db_t;
wire	[17:0]	c1r3_q_t;
wire		c1r3_reg_ena;
wire		c1r3_reg_enb;
wire		c1r3_wea_t;
wire		c1r3_web_t;
wire	[11:0]	c1r2_aa_t;
wire	[11:0]	c1r2_ab_t;
wire		c1r2_cea_t;
wire		c1r2_ceb_t;
wire		c1r2_clka_inv;
wire		c1r2_clka_n;
wire		c1r2_clkb_inv;
wire		c1r2_clkb_n;
wire	[17:0]	c1r2_da_t;
wire	[17:0]	c1r2_db_ecc;
wire	[17:0]	c1r2_db_t;
wire	[17:0]	c1r2_q_t;
wire		c1r2_reg_ena;
wire		c1r2_reg_enb;
wire		c1r2_wea_t;
wire		c1r2_web_t;
wire	[11:0]	c1r1_aa_t;
wire	[11:0]	c1r1_ab_t;
wire		c1r1_cea_t;
wire		c1r1_ceb_t;
wire		c1r1_clka_inv;
wire		c1r1_clka_n;
wire		c1r1_clkb_inv;
wire		c1r1_clkb_n;
wire	[17:0]	c1r1_da_t;
wire	[17:0]	c1r1_db_ecc;
wire	[17:0]	c1r1_db_t;
wire	[17:0]	c1r1_q_t;
wire		c1r1_reg_ena;
wire		c1r1_reg_enb;
wire		c1r1_wea_t;
wire		c1r1_web_t;
wire		clkreg_a;
wire	[63:0]	i_data;
wire	[7:0]	i_parity;
wire		modeax18_4;
wire		modeax18_3;
wire		modeax18_2;
wire		modeax18_1;
wire		modebx18_4;
wire		modebx18_3;
wire		modebx18_2;
wire		modebx18_1;
wire	[63:0]	o_code;
wire	[7:0]	o_parity;
assign c1r1_clka_n = EMB5K_1_PORTA_CKINV ? !c1r1_clka : c1r1_clka;
assign c1r1_clkb_n = EMB5K_1_PORTB_CKINV ? !c1r1_clkb : c1r1_clkb;
assign c1r2_clka_n = EMB5K_2_PORTA_CKINV ? !c1r2_clka : c1r2_clka;
assign c1r2_clkb_n = EMB5K_2_PORTB_CKINV ? !c1r2_clkb : c1r2_clkb;
assign c1r3_clka_n = EMB5K_3_PORTA_CKINV ? !c1r3_clka : c1r3_clka;
assign c1r3_clkb_n = EMB5K_3_PORTB_CKINV ? !c1r3_clkb : c1r3_clkb;
assign c1r4_clka_n = EMB5K_4_PORTA_CKINV ? !c1r4_clka : c1r4_clka;
assign c1r4_clkb_n = EMB5K_4_PORTB_CKINV ? !c1r4_clkb : c1r4_clkb;

wire [71:0] dangling;
supply0_guts G (
	.gnd	(gnd) 
);
supply1_guts V (
	.vcc	(vcc) 
);

//clk_inv u1_clka_inv (
//	.ck_	(c1r1_clka),
//
//	.ck_n	(c1r1_clka_inv) 
//);
//
//gclk_clk_mux u1_cfg_inv_clka (
//	.ck_i0	(c1r1_clka),
//	.ck_i1	(c1r1_clka_inv),
//	.sel	(EMB5K_1_PORTA_CKINV),
//
//	.ck_out	(c1r1_clka_n) 
//);
//
//clk_inv u1_clkb_inv (
//	.ck_	(c1r1_clkb),
//
//	.ck_n	(c1r1_clkb_inv) 
//);
//
//gclk_clk_mux u1_cfg_inv_clkb (
//	.ck_i0	(c1r1_clkb),
//	.ck_i1	(c1r1_clkb_inv),
//	.sel	(EMB5K_1_PORTB_CKINV),
//
//	.ck_out	(c1r1_clkb_n) 
//);
//
//clk_inv u2_clka_inv (
//	.ck_	(c1r2_clka),
//
//	.ck_n	(c1r2_clka_inv) 
//);
//
//gclk_clk_mux u2_cfg_inv_clka (
//	.ck_i0	(c1r2_clka),
//	.ck_i1	(c1r2_clka_inv),
//	.sel	(EMB5K_2_PORTA_CKINV),
//
//	.ck_out	(c1r2_clka_n) 
//);
//
//clk_inv u2_clkb_inv (
//	.ck_	(c1r2_clkb),
//
//	.ck_n	(c1r2_clkb_inv) 
//);
//
//gclk_clk_mux u2_cfg_inv_clkb (
//	.ck_i0	(c1r2_clkb),
//	.ck_i1	(c1r2_clkb_inv),
//	.sel	(EMB5K_2_PORTB_CKINV),
//
//	.ck_out	(c1r2_clkb_n) 
//);
//
//clk_inv u3_clka_inv (
//	.ck_	(c1r3_clka),
//
//	.ck_n	(c1r3_clka_inv) 
//);
//
//gclk_clk_mux u3_cfg_inv_clka (
//	.ck_i0	(c1r3_clka),
//	.ck_i1	(c1r3_clka_inv),
//	.sel	(EMB5K_3_PORTA_CKINV),
//
//	.ck_out	(c1r3_clka_n) 
//);
//
//clk_inv u3_clkb_inv (
//	.ck_	(c1r3_clkb),
//
//	.ck_n	(c1r3_clkb_inv) 
//);
//
//gclk_clk_mux u3_cfg_inv_clkb (
//	.ck_i0	(c1r3_clkb),
//	.ck_i1	(c1r3_clkb_inv),
//	.sel	(EMB5K_3_PORTB_CKINV),
//
//	.ck_out	(c1r3_clkb_n) 
//);
//
//clk_inv u4_clka_inv (
//	.ck_	(c1r4_clka),
//
//	.ck_n	(c1r4_clka_inv) 
//);
//
//gclk_clk_mux u4_cfg_inv_clka (
//	.ck_i0	(c1r4_clka),
//	.ck_i1	(c1r4_clka_inv),
//	.sel	(EMB5K_4_PORTA_CKINV),
//
//	.ck_out	(c1r4_clka_n) 
//);
//
//clk_inv u4_clkb_inv (
//	.ck_	(c1r4_clkb),
//
//	.ck_n	(c1r4_clkb_inv) 
//);
//
//gclk_clk_mux u4_cfg_inv_clkb (
//	.ck_i0	(c1r4_clkb),
//	.ck_i1	(c1r4_clkb_inv),
//	.sel	(EMB5K_4_PORTB_CKINV),
//
//	.ck_out	(c1r4_clkb_n) 
//);

assign c1r1_reg_ena = PEEK_MODE ? peek_en : c1r1_user_ena;
assign c1r1_reg_enb = PEEK_MODE ? peek_en : c1r1_user_enb;
assign c1r2_reg_ena = PEEK_MODE ? peek_en : c1r2_user_ena;
assign c1r2_reg_enb = PEEK_MODE ? peek_en : c1r2_user_enb;
assign c1r3_reg_ena = PEEK_MODE ? peek_en : c1r3_user_ena;
assign c1r3_reg_enb = PEEK_MODE ? peek_en : c1r3_user_enb;
assign c1r4_reg_ena = PEEK_MODE ? peek_en : c1r4_user_ena;
assign c1r4_reg_enb = PEEK_MODE ? peek_en : c1r4_user_enb;

//gclk_clk_mux u1_cfg_ena (
//	.ck_i0	(c1r1_user_ena),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r1_reg_ena) 
//);
//
//gclk_clk_mux u1_cfg_enb (
//	.ck_i0	(c1r1_user_enb),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r1_reg_enb) 
//);
//
//gclk_clk_mux u2_cfg_ena (
//	.ck_i0	(c1r2_user_ena),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r2_reg_ena) 
//);
//
//gclk_clk_mux u2_cfg_enb (
//	.ck_i0	(c1r2_user_enb),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r2_reg_enb) 
//);
//
//gclk_clk_mux u3_cfg_ena (
//	.ck_i0	(c1r3_user_ena),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r3_reg_ena) 
//);
//
//gclk_clk_mux u3_cfg_enb (
//	.ck_i0	(c1r3_user_enb),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r3_reg_enb) 
//);
//
//gclk_clk_mux u4_cfg_ena (
//	.ck_i0	(c1r4_user_ena),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r4_reg_ena) 
//);
//
//gclk_clk_mux u4_cfg_enb (
//	.ck_i0	(c1r4_user_enb),
//	.ck_i1	(peek_en),
//	.sel	(PEEK_MODE),
//
//	.ck_out	(c1r4_reg_enb) 
//);

emb18k_ext u0_emb_ext (
	.a_addr_ext		(a_addr_ext[1:0]),
	.b_addr_ext		(b_addr_ext[1:0]),
	.c1r1_cea_i		(c1r1_cea),
	.c1r1_wea_i		(c1r1_wea),
	.c1r1_ceb_i		(c1r1_ceb),
	.c1r1_web_i		(c1r1_web),
	.c1r2_cea_i		(c1r2_cea),
	.c1r2_wea_i		(c1r2_wea),
	.c1r2_ceb_i		(c1r2_ceb),
	.c1r2_web_i		(c1r2_web),
	.c1r3_cea_i		(c1r3_cea),
	.c1r3_wea_i		(c1r3_wea),
	.c1r3_ceb_i		(c1r3_ceb),
	.c1r3_web_i		(c1r3_web),
	.c1r4_cea_i		(c1r4_cea),
	.c1r4_wea_i		(c1r4_wea),
	.c1r4_ceb_i		(c1r4_ceb),
	.c1r4_web_i		(c1r4_web),
	.c1r1_clka		(c1r1_clka_n),
	.c1r1_clkb		(c1r1_clkb_n),
	.c1r2_clka		(c1r2_clka_n),
	.c1r2_clkb		(c1r2_clkb_n),
	.c1r3_clka		(c1r3_clka_n),
	.c1r3_clkb		(c1r3_clkb_n),
	.c1r4_clka		(c1r4_clka_n),
	.c1r4_clkb		(c1r4_clkb_n),
	.c1r1_rstna		(c1r1_rstna),
	.c1r1_rstnb		(c1r1_rstnb),
	.c1r2_rstna		(c1r2_rstna),
	.c1r2_rstnb		(c1r2_rstnb),
	.c1r3_rstna		(c1r3_rstna),
	.c1r3_rstnb		(c1r3_rstnb),
	.c1r4_rstna		(c1r4_rstna),
	.c1r4_rstnb		(c1r4_rstnb),
	.c1r1_reg_ena		(c1r1_reg_ena),
	.c1r1_reg_enb		(c1r1_reg_enb),
	.c1r2_reg_ena		(c1r2_reg_ena),
	.c1r2_reg_enb		(c1r2_reg_enb),
	.c1r3_reg_ena		(c1r3_reg_ena),
	.c1r3_reg_enb		(c1r3_reg_enb),
	.c1r4_reg_ena		(c1r4_reg_ena),
	.c1r4_reg_enb		(c1r4_reg_enb),
	.gbl_clear_b		(gbl_clear_b),
	.modeax18_1		(modeax18_1),
	.modebx18_1		(modebx18_1),
	.modeax18_2		(modeax18_2),
	.modebx18_2		(modebx18_2),
	.modeax18_3		(modeax18_3),
	.modebx18_3		(modebx18_3),
	.modeax18_4		(modeax18_4),
	.modebx18_4		(modebx18_4),
	.EMB5K_1_MODEA_SEL	(EMB5K_1_MODEA_SEL[3:0]),
	.EMB5K_3_MODEA_SEL	(EMB5K_3_MODEA_SEL[3:0]),
	.EMB5K_1_PORTA_WR_MODE	(EMB5K_1_PORTA_WR_MODE[1:0]),
	.EMB5K_1_PORTB_WR_MODE	(EMB5K_1_PORTB_WR_MODE[1:0]),
	.EMB5K_3_PORTA_WR_MODE	(EMB5K_3_PORTA_WR_MODE[1:0]),
	.EMB5K_3_PORTB_WR_MODE	(EMB5K_3_PORTB_WR_MODE[1:0]),
	.WIDTH_EXT_MODE01	(WIDTH_EXT_MODE01),
	.WIDTH_EXT_MODE23	(WIDTH_EXT_MODE23),
	.DEPTH_EXT_MODE01	(DEPTH_EXT_MODE01),
	.DEPTH_EXT_MODE23	(DEPTH_EXT_MODE23),
	.FIFO_EN		(FIFO_EN),
	.PEEK_MODE		(PEEK_MODE),
	.EXT_18K		(EXT_18K),
	.EMB5K_1_PORTA_REG_OUT	(EMB5K_1_PORTA_REG_OUT),
	.EMB5K_1_PORTB_REG_OUT	(EMB5K_1_PORTB_REG_OUT),
	.EMB5K_2_PORTA_REG_OUT	(EMB5K_2_PORTA_REG_OUT),
	.EMB5K_2_PORTB_REG_OUT	(EMB5K_2_PORTB_REG_OUT),
	.EMB5K_3_PORTA_REG_OUT	(EMB5K_3_PORTA_REG_OUT),
	.EMB5K_3_PORTB_REG_OUT	(EMB5K_3_PORTB_REG_OUT),
	.EMB5K_4_PORTA_REG_OUT	(EMB5K_4_PORTA_REG_OUT),
	.EMB5K_4_PORTB_REG_OUT	(EMB5K_4_PORTB_REG_OUT),
	.rd_mem_n		(rd_mem_n),
	.wr_mem_n		(wr_mem_n),
	.peek_en		(peek_en),
	.peek_rd_en		(peek_rd_en),
	.rptr			(rptr[13:0]),
	.wptr			(wptr[13:0]),
	.c1r1_aa_i		(c1r1_aa[11:0]),
	.c1r1_ab_i		(c1r1_ab[11:0]),
	.c1r2_aa_i		(c1r2_aa[11:0]),
	.c1r2_ab_i		(c1r2_ab[11:0]),
	.c1r3_aa_i		(c1r3_aa[11:0]),
	.c1r3_ab_i		(c1r3_ab[11:0]),
	.c1r4_aa_i		(c1r4_aa[11:0]),
	.c1r4_ab_i		(c1r4_ab[11:0]),
	.c1r1_da_i		(c1r1_da[17:0]),
	.c1r1_db_i		(c1r1_db[17:0]),
	.c1r2_da_i		(c1r2_da[17:0]),
	.c1r2_db_i		(c1r2_db[17:0]),
	.c1r3_da_i		(c1r3_da[17:0]),
	.c1r3_db_i		(c1r3_db[17:0]),
	.c1r4_da_i		(c1r4_da[17:0]),
	.c1r4_db_i		(c1r4_db[17:0]),
	.c1r1_q_i		(c1r1_q_t[17:0]),
	.c1r2_q_i		(c1r2_q_t[17:0]),
	.c1r3_q_i		(c1r3_q_t[17:0]),
	.c1r4_q_i		(c1r4_q_t[17:0]),

	.c1r1_cea		(c1r1_cea_t),
	.c1r1_wea		(c1r1_wea_t),
	.c1r1_ceb		(c1r1_ceb_t),
	.c1r1_web		(c1r1_web_t),
	.c1r2_cea		(c1r2_cea_t),
	.c1r2_wea		(c1r2_wea_t),
	.c1r2_ceb		(c1r2_ceb_t),
	.c1r2_web		(c1r2_web_t),
	.c1r3_cea		(c1r3_cea_t),
	.c1r3_wea		(c1r3_wea_t),
	.c1r3_ceb		(c1r3_ceb_t),
	.c1r3_web		(c1r3_web_t),
	.c1r4_cea		(c1r4_cea_t),
	.c1r4_wea		(c1r4_wea_t),
	.c1r4_ceb		(c1r4_ceb_t),
	.c1r4_web		(c1r4_web_t),
	.c1r1_aa		(c1r1_aa_t[11:0]),
	.c1r1_ab		(c1r1_ab_t[11:0]),
	.c1r2_aa		(c1r2_aa_t[11:0]),
	.c1r2_ab		(c1r2_ab_t[11:0]),
	.c1r3_aa		(c1r3_aa_t[11:0]),
	.c1r3_ab		(c1r3_ab_t[11:0]),
	.c1r4_aa		(c1r4_aa_t[11:0]),
	.c1r4_ab		(c1r4_ab_t[11:0]),
	.c1r1_da		(c1r1_da_t[17:0]),
	.c1r1_db		(c1r1_db_t[17:0]),
	.c1r2_da		(c1r2_da_t[17:0]),
	.c1r2_db		(c1r2_db_t[17:0]),
	.c1r3_da		(c1r3_da_t[17:0]),
	.c1r3_db		(c1r3_db_t[17:0]),
	.c1r4_da		(c1r4_da_t[17:0]),
	.c1r4_db		(c1r4_db_t[17:0]),
	.c1r1_q			(c1r1_q[17:0]),
	.c1r2_q			(c1r2_q[17:0]),
	.c1r3_q			(c1r3_q[17:0]),
	.c1r4_q			(c1r4_q[17:0]),
	.c1r1_no_a		(c1r1_no_a),
	.c1r1_rstna_t		(c1r1_rstna_t) 
);

ecc_enc_wrap u0_ecc_encoder (
	.ECC_ENC_EN	(ECC_ENC_EN),
	.din		({c1r4_db_t[15:0],  c1r3_db_t[15:0],  c1r2_db_t[15:0],  c1r1_db_t[15:0]}),
	.dinp		({c1r4_db_t[17:16], c1r3_db_t[17:16], c1r2_db_t[17:16], c1r1_db_t[17:16]}),
	.eccindberr	(eccindberr),
	.eccinsberr	(eccinsberr),

	.dino		({c1r4_db_ecc[15:0], c1r3_db_ecc[15:0], c1r2_db_ecc[15:0], c1r1_db_ecc[15:0]}),
	.dinpo		({c1r4_db_ecc[17:16], c1r3_db_ecc[17:16], c1r2_db_ecc[17:16], c1r1_db_ecc[17:16]}) 
);

ecc_dec_wrap u0_ecc_decoder (
	.i_data			(i_data[63:0]),
	.i_parity		(i_parity[7:0]),
	.EMB5K_1_PORTA_REG_OUT	(EMB5K_1_PORTA_REG_OUT),
	.DEC_REG_EN		(DEC_REG_EN),
	.ECC_DEC_EN		(ECC_DEC_EN),
	.c1r1_aa		(c1r1_aa_t[11:0]),
	.read_en		(c1r1_no_a),
	.c1r1_rstna		(c1r1_rstna_t),
	.peek_en		(peek_en),
	.FIFO_EN		(FIFO_EN),
	.PEEK_MODE		(PEEK_MODE),
	.peek_rd_en		(peek_rd_en),
	.c1r1_reg_ena		(c1r1_reg_ena),
	.clkreg_a		(clkreg_a),

	.o_code			(o_code[63:0]),
	.o_parity		(o_parity[7:0]),
	.eccoutsberr		(eccoutsberr),
	.eccoutdberr		(eccoutdberr),
	.err_addr		(err_addr[7:0]) 
);

emb5k_core emb5k_core_1 (
	.clka		(c1r1_clka_n),
	.aa		(c1r1_aa_t[11:0]),
	.da		(c1r1_da_t[17:0]),
	.cea		(c1r1_cea_t),
	.wea		(c1r1_wea_t),
	.clkb		(c1r1_clkb_n),
	.ab		(c1r1_ab_t[11:0]),
	.db		(c1r1_db_ecc[17:0]),
	.ceb		(c1r1_ceb_t),
	.web		(c1r1_web_t),
	.MODEA_SEL	(EMB5K_1_MODEA_SEL[3:0]),
	.MODEB_SEL	(EMB5K_1_MODEB_SEL[3:0]),
	.PORTA_WR_MODE	(EMB5K_1_PORTA_WR_MODE[1:0]),
	.PORTB_WR_MODE	(EMB5K_1_PORTB_WR_MODE[1:0]),
	.DEC_REG_EN	(DEC_REG_EN),
	.PORTA_BYPASS	(EMB5K_1_PORTA_BYPASS),
	.PORTB_BYPASS	(EMB5K_1_PORTB_BYPASS),
	.PORTA_CE	(EMB5K_1_PORTA_CE),
	.PORTB_CE	(EMB5K_1_PORTB_CE),
	.PORTA_PROG	(PORTA_PROG[7:0]),
	.PORTB_PROG	(PORTB_PROG[7:0]),
	.gbl_clear_b	(gbl_clear_b),
	.cf_clk		(gnd),
	.ch1en		(gnd),
	.initial_en	(gnd),
	.initial_in	({28{gnd}}),
	.por_a		(vcc),
	.por_b		(vcc),
	.o_code		(o_code[15:0]),
	.o_parity	(o_parity[1:0]),
	.ECC_DEC_EN	(ECC_DEC_EN),

	.q		(c1r1_q_t[17:0]),
	.init_q		(dangling[17:0]),
	.modeax18	(modeax18_1),
	.modebx18	(modebx18_1),
	.clkreg_a	(clkreg_a),
	.i_data		(i_data[15:0]),
	.i_parity	(i_parity[1:0]) 
);

emb5k_core emb5k_core_2 (
	.clka		(c1r2_clka_n),
	.aa		(c1r2_aa_t[11:0]),
	.da		(c1r2_da_t[17:0]),
	.cea		(c1r2_cea_t),
	.wea		(c1r2_wea_t),
	.clkb		(c1r2_clkb_n),
	.ab		(c1r2_ab_t[11:0]),
	.db		(c1r2_db_ecc[17:0]),
	.ceb		(c1r2_ceb_t),
	.web		(c1r2_web_t),
	.MODEA_SEL	(EMB5K_2_MODEA_SEL[3:0]),
	.MODEB_SEL	(EMB5K_2_MODEB_SEL[3:0]),
	.PORTA_WR_MODE	(EMB5K_2_PORTA_WR_MODE[1:0]),
	.PORTB_WR_MODE	(EMB5K_2_PORTB_WR_MODE[1:0]),
	.DEC_REG_EN	(DEC_REG_EN),
	.PORTA_BYPASS	(EMB5K_2_PORTA_BYPASS),
	.PORTB_BYPASS	(EMB5K_2_PORTB_BYPASS),
	.PORTA_CE	(EMB5K_2_PORTA_CE),
	.PORTB_CE	(EMB5K_2_PORTB_CE),
	.PORTA_PROG	(PORTA_PROG[7:0]),
	.PORTB_PROG	(PORTB_PROG[7:0]),
	.gbl_clear_b	(gbl_clear_b),
	.cf_clk		(gnd),
	.ch1en		(gnd),
	.initial_en	(gnd),
	.initial_in	({28{gnd}}),
	.por_a		(vcc),
	.por_b		(vcc),
	.o_code		(o_code[31:16]),
	.o_parity	(o_parity[3:2]),
	.ECC_DEC_EN	(ECC_DEC_EN),

	.q		(c1r2_q_t[17:0]),
	.init_q		(dangling[35:18]),
	.modeax18	(modeax18_2),
	.modebx18	(modebx18_2),
	.clkreg_a	(),
	.i_data		(i_data[31:16]),
	.i_parity	(i_parity[3:2]) 
);

emb5k_core emb5k_core_3 (
	.clka		(c1r3_clka_n),
	.aa		(c1r3_aa_t[11:0]),
	.da		(c1r3_da_t[17:0]),
	.cea		(c1r3_cea_t),
	.wea		(c1r3_wea_t),
	.clkb		(c1r3_clkb_n),
	.ab		(c1r3_ab_t[11:0]),
	.db		(c1r3_db_ecc[17:0]),
	.ceb		(c1r3_ceb_t),
	.web		(c1r3_web_t),
	.MODEA_SEL	(EMB5K_3_MODEA_SEL[3:0]),
	.MODEB_SEL	(EMB5K_3_MODEB_SEL[3:0]),
	.PORTA_WR_MODE	(EMB5K_3_PORTA_WR_MODE[1:0]),
	.PORTB_WR_MODE	(EMB5K_3_PORTB_WR_MODE[1:0]),
	.DEC_REG_EN	(DEC_REG_EN),
	.PORTA_BYPASS	(EMB5K_3_PORTA_BYPASS),
	.PORTB_BYPASS	(EMB5K_3_PORTB_BYPASS),
	.PORTA_CE	(EMB5K_3_PORTA_CE),
	.PORTB_CE	(EMB5K_3_PORTB_CE),
	.PORTA_PROG	(PORTA_PROG[7:0]),
	.PORTB_PROG	(PORTB_PROG[7:0]),
	.gbl_clear_b	(gbl_clear_b),
	.cf_clk		(gnd),
	.ch1en		(gnd),
	.initial_en	(gnd),
	.initial_in	({28{gnd}}),
	.por_a		(vcc),
	.por_b		(vcc),
	.o_code		(o_code[47:32]),
	.o_parity	(o_parity[5:4]),
	.ECC_DEC_EN	(ECC_DEC_EN),

	.q		(c1r3_q_t[17:0]),
	.init_q		(dangling[53:36]),
	.modeax18	(modeax18_3),
	.modebx18	(modebx18_3),
	.clkreg_a	(),
	.i_data		(i_data[47:32]),
	.i_parity	(i_parity[5:4]) 
);

emb5k_core emb5k_core_4 (
	.clka		(c1r4_clka_n),
	.aa		(c1r4_aa_t[11:0]),
	.da		(c1r4_da_t[17:0]),
	.cea		(c1r4_cea_t),
	.wea		(c1r4_wea_t),
	.clkb		(c1r4_clkb_n),
	.ab		(c1r4_ab_t[11:0]),
	.db		(c1r4_db_ecc[17:0]),
	.ceb		(c1r4_ceb_t),
	.web		(c1r4_web_t),
	.MODEA_SEL	(EMB5K_4_MODEA_SEL[3:0]),
	.MODEB_SEL	(EMB5K_4_MODEB_SEL[3:0]),
	.PORTA_WR_MODE	(EMB5K_4_PORTA_WR_MODE[1:0]),
	.PORTB_WR_MODE	(EMB5K_4_PORTB_WR_MODE[1:0]),
	.DEC_REG_EN	(DEC_REG_EN),
	.PORTA_BYPASS	(EMB5K_4_PORTA_BYPASS),
	.PORTB_BYPASS	(EMB5K_4_PORTB_BYPASS),
	.PORTA_CE	(EMB5K_4_PORTA_CE),
	.PORTB_CE	(EMB5K_4_PORTB_CE),
	.PORTA_PROG	(PORTA_PROG[7:0]),
	.PORTB_PROG	(PORTB_PROG[7:0]),
	.gbl_clear_b	(gbl_clear_b),
	.cf_clk		(gnd),
	.ch1en		(gnd),
	.initial_en	(gnd),
	.initial_in	({28{gnd}}),
	.por_a		(vcc),
	.por_b		(vcc),
	.o_code		(o_code[63:48]),
	.o_parity	(o_parity[7:6]),
	.ECC_DEC_EN	(ECC_DEC_EN),

	.q		(c1r4_q_t[17:0]),
	.init_q		(dangling[71:54]),
	.modeax18	(modeax18_4),
	.modebx18	(modebx18_4),
	.clkreg_a	(),
	.i_data		(i_data[63:48]),
	.i_parity	(i_parity[7:6]) 
);


endmodule

// VPERL: GENERATED_END
//
// module: CARRY_SKIP_IN
//
// description: enable the carry input from below cell or not 
// config:      1 bit to select where carry-in from.
//              set 1'b1 when the le is the first stage of adder.
//
//----------------------------------------------------------------------------

module CARRY_SKIP_IN (
	cin,
	
	c0alt,
	c0ripple,
	cskip4,
	cskip8,
	ripple,
	p47,
	p07,
	p03
`ifdef FM_HACK
	,CIN_BELOW
	,ALLOW_SKIP
`endif
);

output	cin;

input	c0alt;
input	c0ripple;
input	cskip4;
input	cskip8;
input	ripple;
input	p47;
input	p07;
input	p03;


`ifdef CS_FORMALPRO_HACK
    wire CIN_BELOW; 
    wire ALLOW_SKIP; 
`else
     `ifdef  SIMULATION
         reg       CIN_BELOW  = 1'b0;
         reg       ALLOW_SKIP = 1'b0;
     `else
		`ifdef FM_HACK
			input	CIN_BELOW;
			input	ALLOW_SKIP;
		`else
			parameter CIN_BELOW  = 1'b0;
         	parameter ALLOW_SKIP = 1'b0;
		`endif
     `endif
`endif
wire    [2:0]    sel ;
wire        p4;

`ifndef CS_SW_SKEL
    assign p4 = !p47 && !p03;
    assign sel = {!p07,p4,!ripple};
    assign cin = ( ALLOW_SKIP == 1'b0 ) 
                ? ( ( CIN_BELOW == 1'b0 ) 
                    ? c0alt 
                    : c0ripple ) 
                : (  ( CIN_BELOW == 1'b0 ) 
                     ? c0alt 
                     : ( sel == 3'b001 )     
                       ? c0ripple  
                       : ( sel == 3'b010 )     
                         ? cskip4 
                         : ( sel == 3'b100 )     
                           ? cskip8 
                           : 1'bx
                  );

    specify
       
    ( c0alt    =>    cin ) = (0,0);                     
    ( c0ripple =>    cin ) = (0,0);                     
    ( cskip4   =>    cin ) = (0,0);                 
    ( cskip8   =>    cin ) = (0,0);       
    ( p07      =>    cin ) = (0,0);                     
    ( p47      =>    cin ) = (0,0);                    
    ( ripple   =>    cin ) = (0,0);                   
    ( p03       =>    cin ) = (0,0);      
            
    endspecify
    
`endif

endmodule
// module: CARRY_SKIP_OUT
//
// description: the carry output logic 
// config:      share 1 bit with CARRY_SKIP_IN to ignore the skip4/8 from below or not 
//              set to 1'b1 when the below carry-in is used.
//
//----------------------------------------------------------------------------

module CARRY_SKIP_OUT (
	r4outb,
	p4outb,
	p8outb,

	plower4,
	p0b,
	p1b,
	p2b,
	p3b
);    

output r4outb;
output p4outb;
output p8outb;

input plower4;
input p0b;
input p1b;
input p2b;
input p3b;

`ifndef CS_SW_SKEL
    wire  p01 ;
    wire  p23 ;

    assign p01 = ~(p0b|p1b);
    assign p23 = ~(p2b|p3b);
    
    assign r4outb =   p01&p23;
    assign p4outb = !(p01&p23);
    assign p8outb = !(p01&p23&plower4);

    specify
       
        ( p0b =>  r4outb ) = (0,0);                     
        ( p1b =>  r4outb ) = (0,0);                     
        ( p2b =>  r4outb ) = (0,0);                 
        ( p3b =>  r4outb ) = (0,0);
        
        
        ( p0b =>  p4outb ) = (0,0);                     
        ( p1b =>  p4outb ) = (0,0);                     
        ( p2b =>  p4outb ) = (0,0);                 
        ( p3b =>  p4outb ) = (0,0);
        
        ( p0b =>  p8outb ) = (0,0);                     
        ( p1b =>  p8outb ) = (0,0);                     
        ( p2b =>  p8outb ) = (0,0);                 
        ( p3b =>  p8outb ) = (0,0);
        ( plower4 =>  p8outb ) = (0,0);
            
    endspecify

`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFG_CLK_GATING
//
// description: clock gating control
//----------------------------------------------------------------------------

module CFG_CLK_GATING (
    clk,
    en,
    clkout
`ifdef FM_HACK
	,cfg_en
`endif
);

input clk;
input en;
output clkout;

`ifdef FM_HACK
	input	cfg_en;
`else
	`ifndef CS_SW_SKEL
		//1: use en, 0: always enable
		parameter cfg_en = 1'b0;
	`endif
`endif

`ifndef CS_SW_SKEL

`ifndef FM_HACK
    wire GSR;
    glbsr inst( .GSR( GSR )) ;

    reg cfg_en_t;
    initial begin
        cfg_en_t = 1;
        #0.1;
        cfg_en_t = 0;
        @(posedge GSR);
        cfg_en_t = cfg_en;
    end
`else
    wire cfg_en_t = cfg_en;
`endif

reg en_latch;
always @(*) begin
    if(cfg_en_t == 0)
        en_latch <= 1;
    else if (clk == 0)
        en_latch <= en;
end

assign clkout = clk & en_latch;
`endif
endmodule

//----------------------------------------------------------------------------
//
// module: CFG_DYN_SWITCH_S2
//
// description: 2 bit wide 2:1 dynamic switch
// config:      2'b00 = output 0 (const)
//				2'b01 = output i0
//				2'b10 = output i1
//				2'b11 = output dynamic switch (fpsel)
//
//----------------------------------------------------------------------------
module CFG_DYN_SWITCH_S2 (
    o,
    i0,
    i1,
    fpsel
`ifdef FM_HACK
	,SEL
`endif
);

input        i0;
input        i1;
input        fpsel;

output        o;

`ifdef CS_FORMALPRO_HACK
   wire [1:0]  SEL;
`else
	`ifdef FM_HACK
		input	[1:0]	SEL;
	`else
		parameter         SEL = 2'b00;
   		parameter         gclk_mux = 0; //0,1,2,3,4,5,6,7
	`endif
`endif

`ifndef FM_HACK
`ifndef CS_SW_SKEL
assign o = 
            (SEL == 2'b00) ? 1'b0 :
            (SEL == 2'b01) ? i0 :
            (SEL == 2'b10) ? i1 :
            (SEL == 2'b11) ? fpsel ? i1 : i0 : 1'bx;       
`endif
`else
//reg gbl_clear_b=1;
//wire GSR;

//initial begin
//    gbl_clear_b = 1'b0;
//    @(posedge GSR);
//    gbl_clear_b = 1'b1;
//end
wire gbl_clear_b=1;

wire ck0 = i0;
wire ck1 = i1;
wire en0b = ~SEL[0];
wire en0  =  SEL[0];
wire en1b = ~SEL[1];
wire en1  =  SEL[1];

reg sel0_reg, sel1_reg;
reg en_ck0, en_ck1;
reg cdone_gate;

wire sel_1p0n =  fpsel & ~en_ck0;
wire sel_0p1n = ~fpsel & ~en_ck1;

always@(posedge ck0 or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        sel0_reg <= 1'b0;
    else
        sel0_reg <= sel_0p1n;
end

always@(negedge ck0 or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        en_ck0 <= 1'b0;
    else
        en_ck0 <= sel0_reg;
end

always@(posedge ck1 or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        sel1_reg <= 1'b0;
    else
        sel1_reg <= sel_1p0n;
end

always@(negedge ck1 or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        en_ck1 <= 1'b0;
    else
        en_ck1 <= sel1_reg;
end

wire enck0 = en0 & (en1 ? en_ck0 : 1'b1);
wire enck1 = en1 & (en0 ? en_ck1 : 1'b1);

wire ck_sel = {enck1, enck0} == 2'b01 ? ck0  :
              {enck1, enck0} == 2'b10 ? ck1  :
              {enck1, enck0} == 2'b00 ? 1'b0 : 1'bx;

always@(negedge ck_sel or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        cdone_gate <= 1'b0;
    else
        cdone_gate <= 1'b1;
end

assign o = cdone_gate & ck_sel;
`endif

endmodule

//----------------------------------------------------------------------------
//
// module: CFGINV
//
// description: configurable inverter
// config:      1 bit to select the invert
//----------------------------------------------------------------------------

module CFGINV (
	o,
	
	i
`ifdef FM_HACK
	,SEL
`endif
);

output	o;

input	i;

`ifdef CS_FORMALPRO_HACK
    wire SEL;
`else
     `ifdef  SIMULATION
          reg       SEL = 1'b1;
     `else
		`ifdef FM_HACK
			input	SEL;
		`else
			parameter SEL = 1'b1;
			parameter         PCK_LOCATION = "NONE";
    		parameter         PLACE_LOCATION = "NONE";
    		parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o = (SEL == 1'b1) ? !i : i;
`endif


endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX10_cmos
//
// description: 1 bit wide 10:1 mux, with additional constant input DEF
// config:      10 bits to select the input (one hot), 
//
//----------------------------------------------------------------------------
module CFGMUX10_cmos (
        o,
        
        i0,
        i1,
        i2,
        i3,
        i4,
        i5,
        i6,
        i7,
        i8,
        i9
`ifdef FM_HACK
        ,SEL
`endif
        );

output        o;

input        i0;
input        i1;
input        i2;
input        i3;
input        i4;
input        i5;
input        i6;
input        i7;
input        i8;
input        i9;

`ifdef CS_FORMALPRO_HACK
    wire [9:0]   SEL;
    wire         DEF;
`else
     `ifdef  SIMULATION
          reg [9:0] SEL = 10'b0000000000;
     `else
        `ifdef FM_HACK
            input    [9:0]    SEL;
        `else
            parameter SEL = 10'b0000000000;
            parameter         CS_PRIM = "bool true";
        `endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign      o   = (SEL == 10'b0000000001) ? i0 :
                      (SEL == 10'b0000000010) ? i1 :
                      (SEL == 10'b0000000100) ? i2 :
                      (SEL == 10'b0000001000) ? i3 : 
                      (SEL == 10'b0000010000) ? i4 :
                      (SEL == 10'b0000100000) ? i5 :
                      (SEL == 10'b0001000000) ? i6 :
                      (SEL == 10'b0010000000) ? i7 :
                      (SEL == 10'b0100000000) ? i8 :
                      (SEL == 10'b1000000000) ? i9 :
                      (SEL == 10'b0000000000) ? 1'bz :                      
                      1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX10S4
//
// description: 1 bit wide 10:1 mux with 4 select
//
//----------------------------------------------------------------------------
module CFGMUX10S4 (
    o,
    i0,
    i1,
    i2,
    i3,
    i4,
    i5,
    i6,
    i7,
    i8,
    i9
`ifdef FM_HACK
	,SEL
`endif
);
   
input i0;
input i1;
input i2;
input i3;
input i4;
input i5;
input i6;
input i7;
input i8;
input i9;

output o;
   
`ifdef CS_FORMALPRO_HACK
    wire [3:0] SEL;
`else
     `ifdef  SIMULATION
          reg [3:0]  SEL = 4'b0000;
     `else
		`ifdef FM_HACK
			input	[3:0]	SEL;
		`else
			parameter  SEL = 4'b0000;
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 4'b0000) ? i0 :
                 (SEL == 4'b0001) ? i1 :
                 (SEL == 4'b0010) ? i2 :
                 (SEL == 4'b0011) ? i3 :
                 (SEL == 4'b0100) ? i4 :
                 (SEL == 4'b0101) ? i5 :
                 (SEL == 4'b0110) ? i6 :
                 (SEL == 4'b0111) ? i7 :
                 (SEL == 4'b1000) ? i8 :
                 (SEL == 4'b1010) ? i8 :
                 (SEL == 4'b1100) ? i8 :
                 (SEL == 4'b1110) ? i8 :
                 (SEL == 4'b1001) ? i9 :
                 (SEL == 4'b1011) ? i9 :
                 (SEL == 4'b1101) ? i9 :
                 (SEL == 4'b1111) ? i9 : 1'bx;
`endif
   
endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX12_43
//
// description: 1 bit wide 6:1 mux, divided into two stages 
// config:      5 bits to select the input, 3 bits 1st stage, 2 bits 2nd stage 
//              (one hot per stage).  
//
//----------------------------------------------------------------------------
module CFGMUX12_43 (
	o,
	i0,
	i1,
	i2,
	i3,
	i4,
	i5,
	i6,
	i7,
	i8,
	i9,
	i10,
	i11
`ifdef FM_HACK
	,SEL
`endif
);

input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11;
output o;
`ifdef CS_FORMALPRO_HACK
   wire [6:0] SEL;
`else
     `ifdef SIMULATION
	  reg [6:0] SEL = 7'b00000;
     `else
		`ifdef FM_HACK
			input [6:0] SEL;
		`else
			parameter SEL = 7'b00000;
		`endif
     `endif
`endif 

`ifndef CS_SW_SKEL
   wire Z0,Z1,Z2;
   assign        Z0 =
                 (SEL[3:0] == 4'b0001) ? i0 :
                 (SEL[3:0] == 4'b0010) ? i1 :
                 (SEL[3:0] == 4'b0100) ? i2 : 
                 (SEL[3:0] == 4'b1000) ? i3 : 
                 (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
   assign        Z1 =
                 (SEL[3:0] == 4'b0001) ? i4 :
                 (SEL[3:0] == 4'b0010) ? i5 :
                 (SEL[3:0] == 4'b0100) ? i6 : 
                 (SEL[3:0] == 4'b1000) ? i7 : 
                 (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
   assign        Z2 =
                 (SEL[3:0] == 4'b0001) ? i8 :
                 (SEL[3:0] == 4'b0010) ? i9 :
                 (SEL[3:0] == 4'b0100) ? i10: 
                 (SEL[3:0] == 4'b1000) ? i11: 
                 (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
   assign	 o =
                 (SEL[6:4] == 3'b001) ? Z0 :
                 (SEL[6:4] == 3'b010) ? Z1 :
                 (SEL[6:4] == 3'b100) ? Z2 :
                 (SEL[6:4] == 3'b000) ? 1'b0 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX16K
//
// description: 1 bit wide 16:1 mux, divided into two stages, with additional
//              input inalt, and constant input DEF.
// config:      9 bits to select the input, 4 bits first stage, 5 bits second
//              stage (one hot per stage).  9'b00000000 selects DEF input, 
//              which is used to source constants. (Should be VCC.)
//              (inalt should be connected to GND.)
//
//----------------------------------------------------------------------------
module CFGMUX16K (
    o,
    i0,
    i1,
    i2,
    i3,
    inalt
`ifdef FM_HACK
	,SEL0
	,SEL1
`endif
);
   
input [3:0]    i0;
input [3:0]     i1;
input [3:0]     i2;
input [3:0]     i3;
input     inalt;

output     o;
   
   // 9 bits per CFGMUX16K
   // 1 x (4 + 4) = 8 CFGMUX16K per ixbar64x32
   // 9 x 8 x 4 = 288 per ixbar
`ifdef CS_FORMALPRO_HACK
    wire [3:0]     SEL0;
    wire [4:0]     SEL1;
    wire         DEF;
`else
     `ifdef  SIMULATION
          reg [3:0] SEL0 = 4'b0000;
          reg [4:0] SEL1 = 5'b00000;
     `else
		`ifdef FM_HACK
			input [3:0] SEL0;
          	input [4:0] SEL1;
		`else
			parameter SEL0 = 4'b0000;
          	parameter SEL1 = 5'b00000;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL
    wire [3:0]     Y;
 
    assign     Y =
           (SEL0 == 4'b0001) ? i0 :
           (SEL0 == 4'b0010) ? i1 :
           (SEL0 == 4'b0100) ? i2 :
           (SEL0 == 4'b1000) ? i3 :
           (SEL0 == 4'b0000) ? 4'b1111 : 4'bxxxx; // dangerous
 
    assign     o =
             (SEL1 == 5'b00001) ? Y[0] :
             (SEL1 == 5'b00010) ? Y[1] :
             (SEL1 == 5'b00100) ? Y[2] :
             (SEL1 == 5'b01000) ? Y[3] :
             (SEL1 == 5'b10000) ? inalt:
             (SEL1 == 5'b00000) ? 1'b1 : 1'bx;
`endif
   
endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX16S4
//
// description: 1 bit wide 16:1 mux
// config:      4 bits to select the input
//
//----------------------------------------------------------------------------
module CFGMUX16S4 (
    o,
    i 
`ifdef FM_HACK
	,SEL
`endif
);
   
input [15:0]    i;
   
output     o;

`ifdef CS_FORMALPRO_HACK
   wire [3:0]     SEL;
   wire         DEF;
`else
     `ifdef  SIMULATION
          reg [3:0] SEL = 4'b0000;
     `else
		`ifdef FM_HACK
			input [3:0] SEL;
		`else
			parameter SEL = 4'b0000;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL   
    assign         o =
                 (SEL == 4'b0000) ? i[0] :
                 (SEL == 4'b0001) ? i[1] :
                 (SEL == 4'b0010) ? i[2] :
                 (SEL == 4'b0011) ? i[3] :
                 (SEL == 4'b0100) ? i[4] :
                 (SEL == 4'b0101) ? i[5] :
                 (SEL == 4'b0110) ? i[6] :
                 (SEL == 4'b0111) ? i[7] :
                 (SEL == 4'b1000) ? i[8] :
                 (SEL == 4'b1001) ? i[9] :
                 (SEL == 4'b1010) ? i[10] :
                 (SEL == 4'b1011) ? i[11] :
                 (SEL == 4'b1100) ? i[12] :
                 (SEL == 4'b1101) ? i[13] :
                 (SEL == 4'b1110) ? i[14] :
                 (SEL == 4'b1111) ? i[15] : 1'bx;
`endif
   
   
endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX16
//
// description: 1 bit wide 16:1 mux, divided into two stages 
// config:      8 bits to select the input, 4 bits per stage 
//              (one hot per stage).  
//
//----------------------------------------------------------------------------
module CFGMUX16 (
    o,
    i0,
    i1,
    i2,
    i3
`ifdef FM_HACK
	,SEL0
	,SEL1
`endif
);
   
input [3:0]    i0;
input [3:0]     i1;
input [3:0]     i2;
input [3:0]     i3;
   
output     o;
   // 8 bits per CFGMUX16
   // 3 x (4 + 4) = 24 CFGMUX16 per ixbar64x32
   // 8 x 24 x 4 = 768 per ixbar
`ifdef CS_FORMALPRO_HACK
   wire [3:0]     SEL0;
   wire [3:0]     SEL1;
   wire         DEF;
`else
     `ifdef  SIMULATION
          reg [3:0] SEL0 = 4'b0000;
          reg [3:0] SEL1 = 4'b0000;
     `else
		`ifdef FM_HACK
			input [3:0] SEL0;
          	input [3:0] SEL1;
		`else
			parameter SEL0 = 4'b0000;
          	parameter SEL1 = 4'b0000;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL   
   wire [3:0]     X;
 
   assign     X =
           (SEL0 == 4'b0001) ? i0 :
           (SEL0 == 4'b0010) ? i1 :
           (SEL0 == 4'b0100) ? i2 :
           (SEL0 == 4'b1000) ? i3 :
           (SEL0 == 4'b0000) ? 4'b1111 : 4'bxxxx; // dangerous
 assign     o =
             (SEL1 == 4'b0001) ? X[0] :
             (SEL1 == 4'b0010) ? X[1] :
             (SEL1 == 4'b0100) ? X[2] :
             (SEL1 == 4'b1000) ? X[3] : 
             (SEL1 == 4'b0000) ? 1'b1 : 1'bx;
`endif
   
   
endmodule
module CFGMUX20I0 (
	in0,
	in1,
	in2,
	in3,
	out
`ifdef FM_HACK
	,SEL0
	,SEL1
`endif
);

output	out;
input	[4:0] in0,in1,in2,in3;
`ifdef FM_HACK
	input [4:0] SEL0;
	input [3:0] SEL1;
`else 
	parameter SEL0 = 5'b00000;
	parameter SEL1 = 4'b0000;
`endif

`ifndef CS_SW_SKEL
wire pg0,pg1,pg2,pg3;

assign 	pg0 = 
	SEL0 == 5'b00001 ? in0[0] :
	SEL0 == 5'b00010 ? in0[1] :
	SEL0 == 5'b00100 ? in0[2] :
	SEL0 == 5'b01000 ? in0[3] :
	SEL0 == 5'b10000 ? in0[4] :
        1'bx;

assign 	pg1 = 
	SEL0 == 5'b00001 ? in1[0] :
	SEL0 == 5'b00010 ? in1[1] :
	SEL0 == 5'b00100 ? in1[2] :
	SEL0 == 5'b01000 ? in1[3] :
	SEL0 == 5'b10000 ? in1[4] :
        1'bx;
assign 	pg2 = 
	SEL0 == 5'b00001 ? in2[0] :
	SEL0 == 5'b00010 ? in2[1] :
	SEL0 == 5'b00100 ? in2[2] :
	SEL0 == 5'b01000 ? in2[3] :
	SEL0 == 5'b10000 ? in2[4] :
        1'bx;
assign 	pg3 = 
	SEL0 == 5'b00001 ? in3[0] :
	SEL0 == 5'b00010 ? in3[1] :
	SEL0 == 5'b00100 ? in3[2] :
	SEL0 == 5'b01000 ? in3[3] :
	SEL0 == 5'b10000 ? in3[4] :
        1'bx;

assign out =
	SEL1 == 4'b0001 ? pg0 :
	SEL1 == 4'b0010 ? pg1 :
	SEL1 == 4'b0100 ? pg2 :
	SEL1 == 4'b1000 ? pg3 :
	SEL1 == 4'b0000 ? 1'b0 :
        1'bx;

`endif
endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX24
//
// description: 1 bit wide 24:1 mux, divided into two stages
// config:      10 bits to select the input, 6 bits first stage, 4 bits second
//              stage (one hot per stage).
//
//----------------------------------------------------------------------------
module CFGMUX24 (
    o,
    i
`ifdef FM_HACK
        ,SEL
`endif
);

input [23:0]  i;
output        o;

 `ifdef CS_FORMALPRO_HACK
     wire [9:0]     SEL;
 `else
     `ifdef  SIMULATION
          reg [9:0] SEL = 10'b000000;
     `else
                `ifdef FM_HACK
                        input        [9:0]        SEL;
                `else
                        parameter SEL = 10'b000000;
                `endif
     `endif
 `endif
 
 `ifndef CS_SW_SKEL
     wire [5:0]     X;
     wire [1:0]     Y;
     
    assign      X[0] =
                   (SEL[3:0] == 4'b0001) ? i[0] :
                   (SEL[3:0] == 4'b0010) ? i[1] :
                   (SEL[3:0] == 4'b0100) ? i[2] :
                   (SEL[3:0] == 4'b1000) ? i[3] :
                   (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
    assign      X[1] =
                   (SEL[3:0] == 4'b0001) ? i[4] :
                   (SEL[3:0] == 4'b0010) ? i[5] :
                   (SEL[3:0] == 4'b0100) ? i[6] :
                   (SEL[3:0] == 4'b1000) ? i[7] :
                   (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
    assign      X[2] =
                   (SEL[3:0] == 4'b0001) ? i[8] :
                   (SEL[3:0] == 4'b0010) ? i[9] :
                   (SEL[3:0] == 4'b0100) ? i[10] :
                   (SEL[3:0] == 4'b1000) ? i[11] :
                   (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
    assign      X[3] =
                   (SEL[3:0] == 4'b0001) ? i[12] :
                   (SEL[3:0] == 4'b0010) ? i[13] :
                   (SEL[3:0] == 4'b0100) ? i[14] :
                   (SEL[3:0] == 4'b1000) ? i[15] :
                   (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
    assign      X[4] =
                   (SEL[3:0] == 4'b0001) ? i[16] :
                   (SEL[3:0] == 4'b0010) ? i[17] :
                   (SEL[3:0] == 4'b0100) ? i[18] :
                   (SEL[3:0] == 4'b1000) ? i[19] :
                   (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
    assign      X[5] =
                   (SEL[3:0] == 4'b0001) ? i[20] :
                   (SEL[3:0] == 4'b0010) ? i[21] :
                   (SEL[3:0] == 4'b0100) ? i[22] :
                   (SEL[3:0] == 4'b1000) ? i[23] :
                   (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;

    assign      Y[0] =
                   (SEL[7:4] == 4'b0001) ? X[0] :
                   (SEL[7:4] == 4'b0010) ? X[1] :
                   (SEL[7:4] == 4'b0100) ? X[2] :
                   (SEL[7:4] == 4'b1000) ? X[3] :
                   (SEL[7:4] == 4'b0000) ? 1'b0 : 1'bx;
    assign      Y[1] =
                   (SEL[5:4] == 2'b01) ? X[4] :
                   (SEL[5:4] == 2'b10) ? X[5] :
                   (SEL[5:4] == 2'b00) ? 1'b0 : 1'bx;

    assign         o =
                   (SEL[9:8] == 2'b01) ? Y[0] :
                   (SEL[9:8] == 2'b10) ? Y[1] :
                   (SEL[9:8] == 2'b00) ? 1'b1 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX2I0
//
// description: 2 bit wide 2:1 mux
// config:      2 bit to select the input
//
//----------------------------------------------------------------------------
module CFGMUX2I0 (
		o,
		
		i0,
		i1
`ifdef FM_HACK
		,SEL
`endif
		);

output		o;

input		i0;
input		i1;
   
`ifdef CS_FORMALPRO_HACK
    wire     [1:0]     SEL;
`else
     `ifdef  SIMULATION
          reg [1:0] SEL = 2'b00;
     `else
		`ifdef FM_HACK
			input	[1:0]	SEL;
		`else
			parameter SEL = 2'b00;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif
 
`ifndef CS_SW_SKEL
    assign         o = 
                    (SEL == 2'b10) ? i1 :
                    (SEL == 2'b01) ? i0 : 
					(SEL == 2'b00) ? 1'b0 : 1'bx;
`endif

endmodule

//----------------------------------------------------------------------------
//
// module: CFGMUX2S1
//
// description: 1 bit wide 2:1 mux
// config:      1 bit to select the input
//
//----------------------------------------------------------------------------
module CFGMUX2S1 (
    o,
    i0,
    i1
`ifdef FM_HACK
	,SEL
`endif
);

input        i0;
input        i1;
output        o;
   
`ifdef CS_FORMALPRO_HACK
    wire         SEL;
`else
     `ifdef  SIMULATION
          reg       SEL = 1'b0;
     `else
		`ifdef FM_HACK
			input	SEL;
		`else
			parameter SEL = 1'b0;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL
    assign         o = SEL ? i1 : i0;

`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX2
//
// description: 2 bit wide 2:1 mux
// config:      2 bit to select the input
//
//----------------------------------------------------------------------------
module CFGMUX2 (
		o,
		
		i0,
		i1
`ifdef FM_HACK
		,SEL
`endif
		);

output		o;

input		i0;
input		i1;
   
`ifdef CS_FORMALPRO_HACK
    wire     [1:0]     SEL;
`else
     `ifdef  SIMULATION
          reg [1:0] SEL = 2'b00;
     `else
		`ifdef FM_HACK
			input	[1:0]	SEL;
		`else
			parameter SEL = 2'b00;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif
 
`ifndef CS_SW_SKEL
    assign         o = 
                    (SEL == 2'b10) ? i1 :
                    (SEL == 2'b01) ? i0 : 
					(SEL == 2'b00) ? 1'b1 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX3I0
//
// description: 1 bit wide 3:1 mux with intial value '0'
// config:      3 bits to select the input (one hot)
//
//----------------------------------------------------------------------------
module CFGMUX3I0 (
    o ,
    
    i0 ,
    i1 ,
    i2
`ifdef FM_HACK
    ,SEL
`endif
);

output    o ;

input    i0 ;
input    i1 ;
input    i2 ;
   
`ifdef CS_FORMALPRO_HACK
    wire [2:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [2:0] SEL = 3'b000;
     `else
        `ifdef FM_HACK
            input    [2:0]    SEL;
        `else
            parameter SEL = 3'b000;
        `endif
     `endif
`endif
 
`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 3'b001) ? i0 :
                 (SEL == 3'b010) ? i1 :
                 (SEL == 3'b100) ? i2 : 
                 (SEL == 3'b000) ? 1'b0 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX3I1
//
// description: 1 bit wide 3:1 mux with intial value '1'
// config:      3 bits to select the input (one hot)
//
//----------------------------------------------------------------------------
module CFGMUX3I1 (
    o ,
    
    i0 ,
    i1 ,
    i2
`ifdef FM_HACK
    ,SEL
`endif
);

output    o ;

input    i0 ;
input    i1 ;
input    i2 ;
   
`ifdef CS_FORMALPRO_HACK
    wire [2:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [2:0] SEL = 3'b000;
     `else
        `ifdef FM_HACK
            input    [2:0]    SEL;
        `else
            parameter SEL = 3'b000;
        `endif
     `endif
`endif
 
`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 3'b001) ? i0 :
                 (SEL == 3'b010) ? i1 :
                 (SEL == 3'b100) ? i2 : 
                 (SEL == 3'b000) ? 1'b1 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX3
//
// description: 1 bit wide 3:1 mux
// config:      3 bits to select the input (one hot)
//
//----------------------------------------------------------------------------
module CFGMUX3 (
	o ,
	
	i0 ,
	i1 ,
	i2
`ifdef FM_HACK
	,SEL
`endif
);

output	o ;

input	i0 ;
input	i1 ;
input	i2 ;
   
`ifdef CS_FORMALPRO_HACK
    wire [2:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [2:0] SEL = 3'b000;
     `else
		`ifdef FM_HACK
			input	[2:0]	SEL;
		`else
			parameter SEL = 3'b000;
		`endif
     `endif
`endif
 
`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 3'b001) ? i0 :
                 (SEL == 3'b010) ? i1 :
                 (SEL == 3'b100) ? i2 : 
                 (SEL == 3'b000) ? 1'b1 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX4_GCO
//
// description: 1 bit wide 4:1 mux, for GCO only
// config:      4 bits to select the input (one hot). 
//
//----------------------------------------------------------------------------
module CFGMUX4_GCO (
		o,

		i0,
		i1,
		i2,
		i3
`ifdef FM_HACK
		,SEL
`endif
		);

output		o;

input		i0;
input		i1;
input		i2;
input		i3;

`ifdef CS_FORMALPRO_HACK
	wire	[3:0]	SEL;
`else
	`ifdef SIMULATION
		reg	[3:0]	SEL = 4'b0000;
	`else
		`ifdef FM_HACK
			input	[3:0]	SEL;
		`else
			parameter SEL = 4'b0000;
		`endif
	`endif
`endif

`ifndef CS_SW_SKEL
wire [1:0] Z;
    assign      Z[0] = 
                    (SEL[1:0] == 2'b10) ? i1 :
                    (SEL[1:0] == 2'b01) ? i0 : 
                    (SEL[1:0] == 2'b00) ? 1'b0 : 1'bx;
    assign      Z[1] = 
                    (SEL[1:0] == 2'b10) ? i3 :
                    (SEL[1:0] == 2'b01) ? i2 : 
                    (SEL[1:0] == 2'b00) ? 1'b0 : 1'bx;

    assign      o    = 
                    (SEL[3:2] == 2'b10) ? Z[1] :
                    (SEL[3:2] == 2'b01) ? Z[0] :
                    (SEL[3:2] == 2'b00) ? 1'b0 : 1'bx;
`endif

endmodule

//----------------------------------------------------------------------------
//
// module: CFGMUX6S5
//
// description: 1 bit wide 4:1 mux with 2 select
// notes:       this is not routing mux
//
//----------------------------------------------------------------------------
module CFGMUX4S2 (
    o,
    i0,
    i1,
    i2,
    i3
`ifdef FM_HACK
	,SEL
`endif
);
   
input i0;
input i1;
input i2;
input i3;
   
output o;
   
`ifdef CS_FORMALPRO_HACK
    wire [1:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [1:0] SEL = 2'b00;
     `else
		`ifdef FM_HACK
			input	[1:0]	SEL;
		`else
			parameter SEL = 2'b00;
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 2'b00) ? i0 :
                 (SEL == 2'b01) ? i1 :
                 (SEL == 2'b10) ? i2 :
                 (SEL == 2'b11) ? i3 : 1'bx;
`endif
   
endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX4
//
// description: 1 bit wide 4:1 mux, 
// config:      4 bits to select the input (one hot). 
//
//----------------------------------------------------------------------------
module CFGMUX4 (
		o,
		
		i0,
		i1,
		i2,
		i3
`ifdef FM_HACK
		,SEL
`endif
		);

output		o;

input		i0;
input		i1;
input		i2;
input		i3;

`ifdef CS_FORMALPRO_HACK
    wire [3:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [3:0] SEL = 4'b0000;
     `else
		`ifdef FM_HACK
			input	[3:0]	SEL;
		`else
			parameter SEL = 4'b0000;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o =
                   (SEL == 4'b0001) ? i0 :
                   (SEL == 4'b0010) ? i1 :
                   (SEL == 4'b0100) ? i2 :
                   (SEL == 4'b1000) ? i3 :
				   (SEL == 4'b0000) ? 1'b1 : 1'bx;
`endif


endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX5
//
// description: 1 bit wide 5:1 mux, with additional constant input DEF
// config:      5 bits to select the input (one hot). 4'b00000 selectes the 
//              DEF input, which is used to source constants.
//
//----------------------------------------------------------------------------
module CFGMUX5 (
    o,
    i0,
    i1,
    i2,
    i3,
    i4
`ifdef FM_HACK
	,SEL
`endif
);

input        i0;
input        i1;
input        i2;
input        i3;
input        i4;

output        o;

`ifdef CS_FORMALPRO_HACK
     wire [4:0]         SEL;
     wire             DEF;
`else
     `ifdef  SIMULATION
          reg [4:0] SEL = 5'b00000;
     `else
		`ifdef FM_HACK
			input	[4:0]	SEL;
		`else
			parameter SEL = 5'b00000;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o =
                   (SEL == 5'b00001) ? i0 :
                   (SEL == 5'b00010) ? i1 :
                   (SEL == 5'b00100) ? i2 :
                   (SEL == 5'b01000) ? i3 :
                   (SEL == 5'b10000) ? i4 : 
				   (SEL == 5'b00000) ? 1'b1 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX6_32
//
// description: 1 bit wide 6:1 mux, divided into two stages 
// config:      5 bits to select the input, 3 bits 1st stage, 2 bits 2nd stage 
//              (one hot per stage).  
//
//----------------------------------------------------------------------------
module CFGMUX6_32 (
	o,
	i0,
	i1,
	i2,
	i3,
	i4,
	i5
`ifdef FM_HACK
	,SEL
`endif
);

input i0,i1,i2,i3,i4,i5;
output o;
`ifdef CS_FORMALPRO_HACK
   wire [4:0] SEL;
`else
     `ifdef SIMULATION
	  reg [4:0] SEL = 5'b00000;
     `else
		`ifdef FM_HACK
			input [4:0] SEL;
		`else
			parameter SEL = 5'b00000;
		`endif
     `endif
`endif 

`ifndef CS_SW_SKEL
   wire Z0,Z1;
   assign        Z0 =
                 (SEL[2:0] == 3'b001) ? i0 :
                 (SEL[2:0] == 3'b010) ? i1 :
                 (SEL[2:0] == 3'b100) ? i2 : 
                 (SEL[2:0] == 3'b000) ? 1'b1 : 1'bx;
   assign        Z1 =
                 (SEL[2:0] == 3'b001) ? i3 :
                 (SEL[2:0] == 3'b010) ? i4 :
                 (SEL[2:0] == 3'b100) ? i5 : 
                 (SEL[2:0] == 3'b000) ? 1'b1 : 1'bx;
   assign	 o =
                 (SEL[4:3] == 2'b01) ? Z0 :
                 (SEL[4:3] == 2'b10) ? Z1 :
                 (SEL[4:3] == 2'b00) ? 1'b0 : 1'bx;
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX6
//
// description: 1 bit wide 6:1 mux, with additional constant input DEF
// config:      6 bits to select the input (one hot), 
//
//----------------------------------------------------------------------------
module CFGMUX6 (
	o,
	
	i0,
	i1,
	i2,
	i3,
	i4,
	i5
`ifdef FM_HACK
	,SEL
`endif
);

output	o;

input	i0;
input	i1;
input	i2;
input	i3;
input	i4;
input	i5;
   
`ifdef CS_FORMALPRO_HACK
    wire [5:0]   SEL;
    wire         DEF;
`else
     `ifdef  SIMULATION
          reg [5:0] SEL = 6'b000000;
     `else
		`ifdef FM_HACK
			input	[5:0]	SEL;
		`else
			parameter SEL = 6'b000000;
			parameter         CS_PRIM = "bool true";
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign      o = (SEL == 6'b000001) ? i0 :
                    (SEL == 6'b000010) ? i1 :
                    (SEL == 6'b000100) ? i2 :
                    (SEL == 6'b001000) ? i3 : 
                    (SEL == 6'b010000) ? i4 :
                    (SEL == 6'b100000) ? i5 :
					(SEL == 6'b000000) ? 1'b1 :
                    1'bx;
   
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: CFGMUX8_42
//
// description: 1 bit wide 6:1 mux, divided into two stages 
// config:      5 bits to select the input, 3 bits 1st stage, 2 bits 2nd stage 
//              (one hot per stage).  
//
//----------------------------------------------------------------------------
module CFGMUX8_42 (
	o,
	i0,
	i1,
	i2,
	i3,
	i4,
	i5,
	i6,
	i7
`ifdef FM_HACK
	,SEL
`endif
);

input i0,i1,i2,i3,i4,i5,i6,i7;
output o;
`ifdef CS_FORMALPRO_HACK
   wire [5:0] SEL;
`else
     `ifdef SIMULATION
	  reg [5:0] SEL = 6'b00000;
     `else
		`ifdef FM_HACK
			input [5:0] SEL;
		`else
			parameter SEL = 6'b00000;
		`endif
     `endif
`endif 

`ifndef CS_SW_SKEL
   wire Z0,Z1;
   assign        Z0 =
                 (SEL[3:0] == 4'b0001) ? i0 :
                 (SEL[3:0] == 4'b0010) ? i1 :
                 (SEL[3:0] == 4'b0100) ? i2 : 
                 (SEL[3:0] == 4'b1000) ? i3 : 
                 (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
   assign        Z1 =
                 (SEL[3:0] == 4'b0001) ? i4 :
                 (SEL[3:0] == 4'b0010) ? i5 :
                 (SEL[3:0] == 4'b0100) ? i6 : 
                 (SEL[3:0] == 4'b1000) ? i7 : 
                 (SEL[3:0] == 4'b0000) ? 1'b1 : 1'bx;
   assign	 o =
                 (SEL[5:4] == 2'b01) ? Z0 :
                 (SEL[5:4] == 2'b10) ? Z1 :
                 (SEL[5:4] == 2'b00) ? 1'b0 : 1'bx;
`endif

endmodule

//----------------------------------------------------------------------------
//
// module: CFGMUX8S3
//
// description: 1 bit wide 8:1 mux with 3 select
//
//----------------------------------------------------------------------------
module CFGMUX8S3 (
    o,
    i0,
    i1,
    i2,
    i3,
    i4,
    i5,
    i6,
    i7
`ifdef FM_HACK
	,SEL
`endif
);
   
input i0;
input i1;
input i2;
input i3;
input i4;
input i5;
input i6;
input i7;
   
output o;
   
`ifdef CS_FORMALPRO_HACK
    wire [2:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [2:0] SEL = 2'b00;
     `else
		`ifdef FM_HACK
			input	[2:0]	SEL;
		`else
			parameter SEL = 3'b000;
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 3'b000) ? i0 :
                 (SEL == 3'b001) ? i1 :
                 (SEL == 3'b010) ? i2 :
                 (SEL == 3'b011) ? i3 :
                 (SEL == 3'b100) ? i4 :
                 (SEL == 3'b101) ? i5 :
                 (SEL == 3'b110) ? i6 :
                 (SEL == 3'b111) ? i7 : 1'bx;
`endif
   
endmodule
//----------------------------------------------------------------------------
//
// module: CFG_NOTINV
//
// description: configurable non-inverter
// config:      1 bit to select the invert
//
//----------------------------------------------------------------------------
module CFG_NOTINV (
    o,
	
    i 
`ifdef FM_HACK
	,SEL
`endif
);

output o;

input  i;

`ifdef CS_FORMALPRO_HACK
    wire SEL;
`else
     `ifdef  SIMULATION
          reg       SEL = 1'b0;
     `else
		`ifdef FM_HACK
			input	SEL;
		`else
			parameter SEL = 1'b0;
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o = (SEL == 1'b1) ? i : !i;
`endif


endmodule
module clk_fb_compensate (
	fclk0_il,
	clkfbin
	`ifdef FM_HACK
	,CFG_FBCLK_EN
	,CFG_FBCLK_INV
	`endif
	);
output	fclk0_il;

input	clkfbin;

`ifdef FM_HACK
input CFG_FBCLK_EN;
input CFG_FBCLK_INV;
`else
parameter CFG_FBCLK_EN = 1'b0;
parameter CFG_FBCLK_INV = 1'b0;
`endif

wire	clk_inv;
xor u0(clk_inv,!clkfbin,CFG_FBCLK_INV);
reg		q_ck;
always @(CFG_FBCLK_EN or clk_inv)
	if(clk_inv == 0) q_ck <= CFG_FBCLK_EN;

wire	feckb;
nand u1(feckb,q_ck,clk_inv);
and u2(fclk0_il,!feckb,CFG_FBCLK_EN);

endmodule

module CVLVDS(
    PAD0,
    PAD1,
    TXD0,
    TXD1,
    TED0,
    TED1,
    RXD0,
    RXD1
`ifdef FM_HACK
,NS_LV_0,NS_LV_1,PDR_0,PDR_1,NDR_0,NDR_1,KEEP_0,KEEP_1,IN_DEL_0,IN_DEL_1,OUT_DEL_0,OUT_DEL_1,
LDR,TERM_DIFF_EN,TD,LVDS_TX_EN,CML_TX_EN,RX_LVDS_EN,RX_DIG_EN_0, 
RX_DIG_EN_1,VPCI_EN_0,VPCI_EN_1,TMDS_TX_EN,LVPECL_TX_EN,CMFB_TX_EN,TERM_CML_EN, 
IN_DEL_EN_0,IN_DEL_EN_1,OUT_DEL_EN_0,OUT_DEL_EN_1
`endif
);

inout  PAD0;
inout  PAD1;
input  TXD0;
input  TXD1;
input  TED0;
input  TED1;
output RXD0;
output RXD1;

supply1 VDDIO, VDDCORE;
supply0 VSSIO, VSSCORE;

`ifdef CS_FORMALPRO_HACK

`else
     `ifdef  SIMULATION
          
     `else
       		`ifdef FM_HACK
		input IN_DEL_EN_0;
		input IN_DEL_EN_1;
		input OUT_DEL_EN_0;
		input OUT_DEL_EN_1;
		input [1:0] NS_LV_0;
		input [1:0] NS_LV_1;         // slew rate control
		input [3:0] PDR_0;
		input [3:0] PDR_1;             // driving strength, P
		input [3:0] NDR_0;
		input [3:0] NDR_1;             // driving strength, N
		input [1:0] KEEP_0;
		input [1:0] KEEP_1;           // pullup,pulldown,bus-keeper
		input [3:0] IN_DEL_0;
		input [3:0] IN_DEL_1;       // input delay
		input [3:0] OUT_DEL_0;
		input [3:0] OUT_DEL_1;     // output delay
		input [2:0] LDR;                     // LVDS driving strength
		
		input TERM_DIFF_EN;                  // LVDS term enable
		input [2:0] TD;                      // LVDS term select
		
		input LVDS_TX_EN;                    // LVDS TX enable
		input CML_TX_EN;                     // CML TX enable
		input RX_LVDS_EN;                    // LVDS RX enable
		input RX_DIG_EN_0;
		input RX_DIG_EN_1;       // LVCMOS RX enable
		input TMDS_TX_EN;
		input LVPECL_TX_EN;
		input CMFB_TX_EN;
		input TERM_CML_EN;
		
		input VPCI_EN_0;
		input VPCI_EN_1;           // PCI diode enable
		//--------------
		`else
		parameter IN_DEL_EN_0 = 1'b0;
		parameter IN_DEL_EN_1 = 1'b0;
		parameter OUT_DEL_EN_0 = 1'b0;
		parameter OUT_DEL_EN_1 = 1'b0;
		parameter [1:0] NS_LV_0 = 2'b0;
		parameter [1:0] NS_LV_1 = 2'b0;         // slew rate control
		parameter [3:0] PDR_0 = 4'b0;
		parameter [3:0] PDR_1 = 4'b0;             // driving strength, P
		parameter [3:0] NDR_0 = 4'b0;
		parameter [3:0] NDR_1 = 4'b0;             // driving strength, N
		parameter [1:0] KEEP_0 = 2'b0;
		parameter [1:0] KEEP_1 = 2'b0;           // pullup,pulldown,bus-keeper
		parameter [3:0] IN_DEL_0 = 4'b0;
		parameter [3:0] IN_DEL_1 = 4'b0;       // input delay
		parameter [3:0] OUT_DEL_0 = 4'b0;
		parameter [3:0] OUT_DEL_1 = 4'b0;     // output delay
		parameter [2:0] LDR = 3'b0;                     // LVDS driving strength
		parameter TERM_DIFF_EN = 1'b0;                  // LVDS term enable
		parameter [2:0] TD = 3'b0;                      // LVDS term select
		parameter LVDS_TX_EN = 1'b0;                    // LVDS TX enable
		parameter CML_TX_EN = 1'b0;                     // CML TX enable
		parameter RX_LVDS_EN = 1'b0;                    // LVDS RX enable
		parameter RX_DIG_EN_0 = 1'b0;
		parameter RX_DIG_EN_1 = 1'b0;       // LVCMOS RX enable
		parameter TMDS_TX_EN = 1'b0;
		parameter LVPECL_TX_EN = 1'b0;
		parameter CMFB_TX_EN = 1'b0;
		parameter TERM_CML_EN = 1'b0;
		parameter VPCI_EN_0 = 1'b0;
		parameter VPCI_EN_1 = 1'b0;           // PCI diode enable
		`endif	 	   
     `endif
`endif
 
`ifndef CS_SW_SKEL
    wire rxe0,rxe1;
    
    assign rxe0=~(RX_DIG_EN_0|RX_LVDS_EN);
    bufif1 rx00 (RXD0,PAD0,RX_DIG_EN_0);
    bufif1 rx02 (RXD0,PAD0,RX_LVDS_EN);
    nmos  NMOSrx0 (RXD0, VSSIO, rxe0);

    assign rxe1=~(RX_DIG_EN_1|RX_LVDS_EN);
    bufif1 rx10 (RXD1,PAD1,RX_DIG_EN_1);
    bufif1 rx12 (RXD1,PAD0,RX_LVDS_EN);
    nmos  NMOSrx1 (RXD1, VSSIO, rxe1);


    //--------- term 
    wire terml,termp0,termp1,termn0,termn1;
    
    assign terml=TERM_DIFF_EN;


    rnmos    TNMOS2A    (PAD1,       TPAD2A_out, terml);
    rnmos    TNMOS2B    (TPAD2A_out, TPAD2B_out, terml);
    rnmos    TNMOS2C    (TPAD2B_out, PAD0,       terml);


    //------- driver 
//------LVCMOS  
    wire pdr0a,ndr0a,pdr0b,ndr0b,pdr0c,ndr0c,pdr1a,ndr1a,pdr1b,ndr1b,pdr1c,ndr1c;
      
    assign pdr0a=PDR_0[0]|PDR_0[1]|PDR_0[2]|PDR_0[3];
    assign ndr0a=NDR_0[0]|NDR_0[1]|NDR_0[2]|NDR_0[3];
    assign pdr0b=pdr0a&(NS_LV_0[0]|NS_LV_0[1])&(!TED0);
    assign ndr0b=ndr0a&(NS_LV_0[0]|NS_LV_0[1])&(!TED0);
    assign pdr0c=~( pdr0b & TXD0 );
    assign ndr0c=~(!ndr0b | TXD0 );
    
    pmos  pdriver00 (PAD0, VDDIO, pdr0c);
    nmos  ndriver00 (PAD0, VSSIO, ndr0c);

    assign pdr1a=PDR_1[0]|PDR_1[1]|PDR_1[2]|PDR_1[3];
    assign ndr1a=NDR_1[0]|NDR_1[1]|NDR_1[2]|NDR_1[3];
    assign pdr1b=pdr1a&(NS_LV_1[0]|NS_LV_1[1])&(!TED1);
    assign ndr1b=ndr1a&(NS_LV_1[0]|NS_LV_1[1])&(!TED1);
    assign pdr1c=~( pdr1b & TXD1 );
    assign ndr1c=~(!ndr1b | TXD1 );
    
    pmos  pdriver10 (PAD1, VDDIO, pdr1c);
    nmos  ndriver10 (PAD1, VSSIO, ndr1c);

//------LVDS
    wire ldr,lpdrp0,lpdrp1,lpdrn0,lpdrn1;    
    
    assign ldr=(|LDR)&TED0&(LVDS_TX_EN|CML_TX_EN);
    assign lpdrp0=~(TXD0&ldr);
    assign lpdrn0=~(TXD0|(~ldr));
    assign lpdrp1=~(!TXD0&ldr);
    assign lpdrn1=~(!TXD0|(~ldr));
    

    pmos  pdriverl0 (PAD0, VDDIO, lpdrp0);
    nmos  ndriverl0 (PAD0, VSSIO, lpdrn0);
    pmos  pdriverl1 (PAD1, VDDIO, lpdrp1);
    nmos  ndriverl1 (PAD1, VSSIO, lpdrn1);

    
    //--------- Pullup 
    wire pullup0,pullup1,pulldn0,pulldn1;
    
    assign pullup0=~(KEEP_0[1]&((!KEEP_0[0])|(KEEP_0[0]&!RXD0)));
    assign pullup1=~(KEEP_1[1]&((!KEEP_1[0])|(KEEP_1[0]&!RXD1)));
    
    rpmos    PMOS0A    (PAD0,       PAD0PA_out, pullup0);
    rpmos    PMOS0B    (PAD0PA_out, PAD0PB_out, pullup0);
    rpmos    PMOS0C    (PAD0PB_out, VDDIO,      pullup0);    

    rpmos    PMOS1A    (PAD1,       PAD1PA_out, pullup1);
    rpmos    PMOS1B    (PAD1PA_out, PAD1PB_out, pullup1);
    rpmos    PMOS1C    (PAD1PB_out, VDDIO,      pullup1);    


    //---------- Pulldown (Strength to Weak)
    assign pulldn0=(KEEP_0[0]&((!KEEP_0[1])|(KEEP_0[1]&RXD0)));
    assign pulldn1=(KEEP_1[0]&((!KEEP_1[1])|(KEEP_1[1]&RXD1)));
    
    rnmos    NMOS0A    (PAD0,       PAD0NA_out, pulldn0);
    rnmos    NMOS0B    (PAD0NA_out, PAD0NB_out, pulldn0);
    rnmos    NMOS0C    (PAD0NB_out, VSSIO,      pulldn0);

    rnmos    NMOS1A    (PAD1,       PAD1NA_out, pulldn1);
    rnmos    NMOS1B    (PAD1NA_out, PAD1NB_out, pulldn1);
    rnmos    NMOS1C    (PAD1NB_out, VSSIO,      pulldn1);
`endif


endmodule

//----------------------------------------------------------------------------
//
// module: DIV
//
// description: Logic divider with asynchronous clear input
// config:      TBD
//
//----------------------------------------------------------------------------
module DIV (
    CKOUT,
    CKIN,
    CLR
`ifdef FM_HACK
    ,DIV
`endif
);

output CKOUT;
input  CKIN;
input  CLR;

`ifdef FM_HACK
    input [3:0]  DIV;
`else
    parameter DIV = 4'b0000;
`endif

//function description 
/* ------------
CLR: 1 rst;
DIV: 0000: bypass
     0001: div 1
     0010: div 2
     0011: div 3
     0100: div4
     0101: div5
     0110: div6
     0111: div7
     1000: div8
     1001: div9
     1010: div10
     1011: div11
     1100: div12
     1101: div13
     1110: div14
     1111: div15
------------ */
wire Q1, Q2, Q3, Q4;
wire Q1N, Q2N, Q3N, Q4N;
wire CKOUT1;
wire CKOUT1B;

wire CKOUT = DIV[3:0]==0 ? CKIN : CKOUT1;

wire SET_DIV = (DIV[0] ^ Q1N) & (DIV[1] ^ Q2N) & (DIV[2] ^ Q3N) & (DIV[3] ^ Q4N);
wire net0342 = ~(DIV[0] & CKIN);
wire net0157 = (Q3N ^ DIV[3]) & (Q2N ^ DIV[2]) & (Q1N ^ DIV[1]) & (CKOUT1B ^ 1'b1);

wire SET_DUTY = net0342 & net0157;
wire SET_DIV_DLY = ~CLR & ~SET_DIV;

wire d1 = ~CLR ^ Q1;
wire d2 = (SET_DIV_DLY & Q1) ^ Q2;
wire d3 = (SET_DIV_DLY & Q1 & Q2) ^ Q3;
wire d4 = (SET_DIV_DLY & Q1 & Q2 & Q3) ^ Q4;

cts_dffrs I119 ( .RSTN(SET_DIV_DLY), .SETN(vcc), .CK(CKIN), .D(d1), .QB(Q1N), .Q(Q1));
cts_dffrs I136 ( .RSTN(SET_DIV_DLY), .SETN(vcc), .CK(CKIN), .D(d2), .QB(Q2N), .Q(Q2));
cts_dffrs I137 ( .RSTN(SET_DIV_DLY), .SETN(vcc), .CK(CKIN), .D(d3), .QB(Q3N), .Q(Q3));
cts_dffrs I138 ( .RSTN(SET_DIV_DLY), .SETN(vcc), .CK(CKIN), .D(d4), .QB(Q4N), .Q(Q4));

cts_dffrs I116 ( .RSTN(~CLR), .SETN(~SET_DIV), .CK(SET_DUTY), .D(1'b0), .QB(CKOUT1B), .Q(CKOUT1));

supply1_guts V ( .vcc	(vcc) );


endmodule
// VPERL: GENERATED_BEG

module DLLV1(
	DLL_CKOUT1,
	DLL_CKOUT0,
	DLLCK,
	DQS
`ifdef FM_HACK
    ,MDLL_BK
    ,MDLL_DR
    ,MDLL_DTEST_EN
    ,MDLL_DTEST_SEL
    ,MDLL_FBSEL
    ,MDLL_MSEL
    ,MDLL_START
    ,SDLL_BK
    ,SDLL_DOFF
    ,SDLL_SSEL
    ,SDLL_START_S
    ,MDLL_MUX_SEL
`endif
);

output		DLL_CKOUT1;
output		DLL_CKOUT0;
input		DLLCK;
input		DQS;
`ifdef FM_HACK
input [3:0]     MDLL_BK;
input           MDLL_DR;
input           MDLL_DTEST_EN;
input [1:0]     MDLL_DTEST_SEL;
input [1:0]     MDLL_FBSEL;
input [3:0]     MDLL_MSEL;
input           MDLL_START;
input [1:0]     SDLL_BK;
input [4:0]     SDLL_DOFF;
input [3:0]     SDLL_SSEL;
input           SDLL_START_S;
input [1:0]     MDLL_MUX_SEL;
`else
parameter      MDLL_BK           = 4'b0 ;
parameter      MDLL_DR           = 1'b0 ;
parameter      MDLL_DTEST_EN     = 1'b0 ;
parameter      MDLL_DTEST_SEL    = 2'b0 ;
parameter      MDLL_FBSEL        = 2'b0 ;
parameter      MDLL_MSEL         = 4'b0 ;
parameter      MDLL_START        = 1'b0 ;
parameter      SDLL_BK           = 2'b0 ;
parameter      SDLL_DOFF         = 5'b0 ;
parameter      SDLL_SSEL         = 4'b0 ;
parameter      SDLL_START_S      = 1'b0 ;
parameter      MDLL_MUX_SEL      = 2'b0 ;
`endif
wire	[18:0]	dangling;

MDLLV1 MDLL (
	.DLLCK		(DLLCK),
	.BK		(MDLL_BK[3:0]),
	.DR		(MDLL_DR),
	.DTEST_EN	(MDLL_DTEST_EN),
	.DTEST_SEL	(MDLL_DTEST_SEL[1:0]),
	.FBSEL		(MDLL_FBSEL[1:0]),
	.MSEL		(MDLL_MSEL[3:0]),
	.START		(MDLL_START),

	.CKOUT		(DLL_CKOUT0),
	.CLKUP		(dangling[5]),
	.DCTLO		(dangling[15:6]),
	.DLOCK		(dangling[4]),
	.DTEST		(dangling[16]),
	.FAIL		(dangling[3]),
	.OF		(dangling[17]),
	.UF		(dangling[18]) 
);

SDLLV1 SDLL (
	.CLKUP		(dangling[5]),
	.DCTLIN		(dangling[15:6]),
	.DQS		(DQS),
	.BK		(SDLL_BK[1:0]),
	.DOFF		(SDLL_DOFF[4:0]),
	.FBSEL		(MDLL_FBSEL[1:0]),
	.SSEL		(SDLL_SSEL[3:0]),
	.START_S	(SDLL_START_S),

	.DQS_O		(DLL_CKOUT1),
	.SOF		(dangling[2]),
	.SUF		(dangling[1]) 
);

endmodule

// VPERL: GENERATED_END
//DSP arch model for QC family
// 20140616: remove underscore in portname, imctrl[4:0]=>imctrl[5:0]

module DSP56V1 (
	alcasout,
	aucasout,
	clcasout,
	cucasout,
	imatch,
	match,
	overflow,
	r,
	rcarrycasout,
	rcasout,
	recarrycasout,
	underflow,
	al,
	alcasin,
	au,
	aucasin,
	cecomp,
	ceibuf,
	cemultl,
	cemultu,
	cepoa,
	cepra,
	ceufc,
	cl,
	clcasin,
	clk,
	cu,
	cucasin,
	dl,
	du,
	ialuctrl,
	iblctrl,
	ibuctrl,
	icctrl,
	ifcctrl,
	ifrctrl,
	imctrl,
	iparctrl,
	ipasctrl,
	ipasubctrl,
	ipazctrl,
	irndm,
	isubctrl,
	iufcctrl,
	rcarrycasin,
	rcasin,
	recarrycasin,
	rstn,
	u 
`ifdef FM_HACK
    ,cfg_pra_au
    ,cfg_pra_cu
    ,cfg_pra_du
    ,cfg_pra_dl
    ,cfg_pra_al
    ,cfg_pra_cl
    ,cfg_pra_ou
    ,cfg_pra_ol
    ,cfg_mult_u
    ,cfg_mult_l
    ,cfg_ufcmux
    ,cfg_vldbit
    ,cfg_match
    ,cfg_imatch
    ,cfg_poa_cyout
    ,cfg_poa_rout
    ,cfg_poa_ceyout
    ,cfg_poa_ceyin
    ,cfg_mat_clr
    ,cfg_pazctrl
    ,cfg_parctrl
    ,cfg_pasubctrl
    ,cfg_blctrl
    ,cfg_buctrl
    ,cfg_pasctrl
    ,cfg_aluctrl
    ,cfg_fcctrl
    ,cfg_ufcctrl
    ,cfg_subctrl
    ,cfg_mctrl
    ,cfg_cctrl
    ,cfg_frctrl
    ,cfg_rndm
`endif
);

output	[17:0]	alcasout;
output	[17:0]	aucasout;
output	[17:0]	clcasout;
output	[17:0]	cucasout;
output		imatch;
output		match;
output		overflow;
output	[71:0]	r;
output		rcarrycasout;
output	[55:0]	rcasout;
output		recarrycasout;
output		underflow;
input	[17:0]	al;
input	[17:0]	alcasin;
input	[17:0]	au;
input	[17:0]	aucasin;
input		cecomp;
input		ceibuf;
input		cemultl;
input		cemultu;
input		cepoa;
input		cepra;
input		ceufc;
input	[17:0]	cl;
input	[17:0]	clcasin;
input		clk;
input	[17:0]	cu;
input	[17:0]	cucasin;
input	[17:0]	dl;
input	[17:0]	du;
input	[2:0]	ialuctrl;
input		iblctrl;
input		ibuctrl;
input	[2:0]	icctrl;
input	[2:0]	ifcctrl;
input	[1:0]	ifrctrl;
input	[5:0]	imctrl;
input	[5:0]	iparctrl;
input	[7:0]	ipasctrl;
input	[1:0]	ipasubctrl;
input	[5:0]	ipazctrl;
input		irndm;
input	[2:0]	isubctrl;
input		iufcctrl;
input		rcarrycasin;
input	[55:0]	rcasin;
input		recarrycasin;
input		rstn;
input	[55:0]	u;

`ifdef FM_HACK
    input [2:0]    cfg_pra_au     ;
    input [2:0]    cfg_pra_cu     ;
    input          cfg_pra_du     ;
    input          cfg_pra_dl     ;
    input [2:0]    cfg_pra_al     ;
    input [2:0]    cfg_pra_cl     ;
    input          cfg_pra_ou     ;
    input          cfg_pra_ol     ;
    input [1:0]    cfg_mult_u     ;
    input [1:0]    cfg_mult_l     ;
    input          cfg_ufcmux     ;
    input [55:0]    cfg_vldbit     ;
    input          cfg_match      ;
    input          cfg_imatch     ;
    input          cfg_poa_cyout  ;
    input [1:0]    cfg_poa_rout   ;
    input          cfg_poa_ceyout ;
    input          cfg_poa_ceyin  ;
    input          cfg_mat_clr    ;
    input          cfg_pazctrl    ;
    input          cfg_parctrl    ;
    input          cfg_pasubctrl  ;
    input          cfg_blctrl     ;
    input          cfg_buctrl     ;
    input          cfg_pasctrl    ;
    input          cfg_aluctrl    ;
    input          cfg_fcctrl     ;
    input          cfg_ufcctrl    ;
    input          cfg_subctrl    ;
    input          cfg_mctrl      ;
    input          cfg_cctrl      ;
    input          cfg_frctrl     ;
    input          cfg_rndm       ;
`else
parameter   cfg_pra_au     = 3'b0;
parameter   cfg_pra_cu     = 3'b0;
parameter   cfg_pra_du     = 1'b0;
parameter   cfg_pra_dl     = 1'b0;
parameter   cfg_pra_al     = 3'b0;
parameter   cfg_pra_cl     = 3'b0;
parameter   cfg_pra_ou     = 1'b0;
parameter   cfg_pra_ol     = 1'b0;
parameter   cfg_mult_u     = 2'b0;
parameter   cfg_mult_l     = 2'b0;
parameter   cfg_ufcmux     = 1'b0;
parameter   cfg_vldbit     = 56'b0;
parameter   cfg_match      = 1'b0;
parameter   cfg_imatch     = 1'b0;
parameter   cfg_poa_cyout  = 1'b0;
parameter   cfg_poa_rout   = 2'b0;
parameter   cfg_poa_ceyout = 1'b0;
parameter   cfg_poa_ceyin  = 1'b0;
parameter   cfg_mat_clr    = 1'b0;
parameter   cfg_pazctrl    = 1'b0;
parameter   cfg_parctrl    = 1'b0;
parameter   cfg_pasubctrl  = 1'b0;
parameter   cfg_blctrl     = 1'b0;
parameter   cfg_buctrl     = 1'b0;
parameter   cfg_pasctrl    = 1'b0;
parameter   cfg_aluctrl    = 1'b0;
parameter   cfg_fcctrl     = 1'b0;
parameter   cfg_ufcctrl    = 1'b0;
parameter   cfg_subctrl    = 1'b0;
parameter   cfg_mctrl      = 1'b0;
parameter   cfg_cctrl      = 1'b0;
parameter   cfg_frctrl     = 1'b0;
parameter   cfg_rndm       = 1'b0;
`endif

dsp_core dsp_core (
	.al		(al[17:0]),
	.alcasin	(alcasin[17:0]),
	.au		(au[17:0]),
	.aucasin	(aucasin[17:0]),
	.cecomp		(cecomp),
	.ceibuf		(ceibuf),
	.cemultl	(cemultl),
	.cemultu	(cemultu),
	.cepoa		(cepoa),
	.cepra		(cepra),
	.ceufc		(ceufc),
	.cfg_aluctrl	(cfg_aluctrl),
	.cfg_blctrl	(cfg_blctrl),
	.cfg_buctrl	(cfg_buctrl),
	.cfg_cctrl	(cfg_cctrl),
	.cfg_fcctrl	(cfg_fcctrl),
	.cfg_frctrl	(cfg_frctrl),
	.cfg_imatch	(cfg_imatch),
	.cfg_mat_clr	(cfg_mat_clr),
	.cfg_match	(cfg_match),
	.cfg_mctrl	(cfg_mctrl),
	.cfg_mult_l	(cfg_mult_l[1:0]),
	.cfg_mult_u	(cfg_mult_u[1:0]),
	.cfg_parctrl	(cfg_parctrl),
	.cfg_pasctrl	(cfg_pasctrl),
	.cfg_pasubctrl	(cfg_pasubctrl),
	.cfg_pazctrl	(cfg_pazctrl),
	.cfg_poa_ceyin	(cfg_poa_ceyin),
	.cfg_poa_ceyout	(cfg_poa_ceyout),
	.cfg_poa_cyout	(cfg_poa_cyout),
	.cfg_poa_rout	(cfg_poa_rout[1:0]),
	.cfg_pra_al	(cfg_pra_al[2:0]),
	.cfg_pra_au	(cfg_pra_au[2:0]),
	.cfg_pra_cl	(cfg_pra_cl[2:0]),
	.cfg_pra_cu	(cfg_pra_cu[2:0]),
	.cfg_pra_dl	(cfg_pra_dl),
	.cfg_pra_du	(cfg_pra_du),
	.cfg_pra_ol	(cfg_pra_ol),
	.cfg_pra_ou	(cfg_pra_ou),
	.cfg_rndm	(cfg_rndm),
	.cfg_subctrl	(cfg_subctrl),
	.cfg_ufcctrl	(cfg_ufcctrl),
	.cfg_ufcmux	(cfg_ufcmux),
	.cfg_vldbit	(cfg_vldbit[55:0]),
	.cl		(cl[17:0]),
	.clcasin	(clcasin[17:0]),
	.clk		(clk),
	.cu		(cu[17:0]),
	.cucasin	(cucasin[17:0]),
	.dl		(dl[17:0]),
	.du		(du[17:0]),
	.ialuctrl	(ialuctrl[2:0]),
	.iblctrl	(iblctrl),
	.ibuctrl	(ibuctrl),
	.icctrl		(icctrl[2:0]),
	.ifcctrl	(ifcctrl[2:0]),
	.ifrctrl	(ifrctrl[1:0]),
	.imctrl		(imctrl[5:0]),
	.iparctrl	(iparctrl[5:0]),
	.ipasctrl	(ipasctrl[7:0]),
	.ipasubctrl	(ipasubctrl[1:0]),
	.ipazctrl	(ipazctrl[5:0]),
	.irndm		(irndm),
	.isubctrl	(isubctrl[2:0]),
	.iufcctrl	(iufcctrl),
	.rcarrycasin	(rcarrycasin),
	.rcasin		(rcasin[55:0]),
	.recarrycasin	(recarrycasin),
	.rstn		(rstn),
	.sck		(gnd),
	.sen		(gnd),
	.si		(gnd),
	.smode		(gnd),
	.srst		(gnd),
	.u		(u[55:0]),

	.alcasout	(alcasout[17:0]),
	.aucasout	(aucasout[17:0]),
	.clcasout	(clcasout[17:0]),
	.cucasout	(cucasout[17:0]),
	.imatch		(imatch),
	.match		(match),
	.overflow	(overflow),
	.r		(r[71:0]),
	.rcarrycasout	(rcarrycasout),
	.rcasout	(rcasout[55:0]),
	.recarrycasout	(recarrycasout),
	.underflow	(underflow) 
);

supply0_guts G (
	.gnd	(gnd) 
);
endmodule


//----------------------------------------------------------------------------
//
// module: efuse_idx16
//
// description: efuse output connecting to FP
//
//----------------------------------------------------------------------------
module efuse_idx16 (
    o 
);

output [15:0]  o;

`ifdef CS_FORMALPRO_HACK
   wire [15:0] 		DATA;
`else
   parameter 	DATA = 16'h0000;
`endif
   
`ifndef CS_SW_SKEL
   assign 		o = DATA;
`endif
   

endmodule
//----------------------------------------------------------------------------
//
// module: EMBMUX5S4
//
// description: 1 bit wide 4:1 mux with 4 select
// notes:       this is not routing mux
//
//----------------------------------------------------------------------------
module EMBMUX5S4 (
    o,  
    i0,  
    i1,  
    i2,  
    i3,  
    i4
`ifdef FM_HACK
		,SEL
`endif
);    
   
input i0;
input i1;
input i2;
input i3;
input i4;

output o;
   
`ifdef CS_FORMALPRO_HACK
    wire     [3:0]     SEL;
`else
     `ifdef  SIMULATION
          reg [3:0] SEL = 4'b0000;
     `else
		`ifdef FM_HACK
			input	[3:0]	SEL;
		`else
			parameter SEL = 4'b0000;
		`endif
     `endif
`endif
   
`ifndef CS_SW_SKEL
   assign               o = 
                             (SEL == 4'b0000) ? i0 : 
                             (SEL == 4'b1000) ? i1 : 
                             (SEL == 4'b1100) ? i2 : 
                             (SEL == 4'b1110) ? i3 : 
                             (SEL == 4'b1111) ? i4 : i4; 
`endif
   
endmodule

//----------------------------------------------------------------------------
//
// module: FG6X2
//
// description: 6 input lookup-table
//        outputs include one of two LUT5 results
// config:      64 bit init value for two LUT5 and 1 bit to select LUT6
//
//----------------------------------------------------------------------------
module FG6X2 (
    x,
    xy,
    f
`ifdef FM_HACK
    ,config_data
    ,mode
`endif
);

    input    [5:0]    f;

    output        x;
    output        xy;


`ifdef CS_FORMALPRO_HACK
    wire [63:0]     config_data;
    wire            mode;
`else
     `ifdef  SIMULATION
          reg [63:0] config_data = 64'h0000000000000000; // [31:0] for LUT5_0, [63:32] for LUT5_1
          reg        mode        = 1'b0;                 // select between LUT6 and LUT5_2
     `else
        `ifdef FM_HACK
            input    [63:0]    config_data;
            input            mode;
        `else
            parameter  [63:0] config_data = 64'h0000000000000000; // [31:0] for LUT5_0, [63:32] for LUT5_1
            parameter  mode        = 1'b0;                 // select between LUT6 and LUT5_2
        `endif
     `endif
`endif

`ifdef SIMULATION    
    reg [63:0] cfg_data;
    initial #1 cfg_data = ~config_data;
`else 
    `ifndef FM_HACK
        localparam [63:0] cfg_data = ~config_data;
    `else
        wire [63:0] cfg_data = ~config_data;
    `endif
`endif

    wire    x0, x1;
    wire        y;

`ifndef CS_SW_SKEL

    
LUT5    lut_0 (
    .f4    (f[4]),
    .f3    (f[3]),
    .f2    (f[2]),
    .f1    (f[1]),
    .f0    (f[0]),
    .dx    (x0)
`ifdef FM_HACK
    ,.config_data (cfg_data[31:0])
`endif
);
`ifndef CS_FORMALPRO_HACK 
     `ifdef  SIMULATION
//        initial  lut_0.config_data=config_data[31:0];
     `else
        `ifdef FM_HACK
        //BLANK param
        `else
            defparam lut_0.config_data=cfg_data[31:0];
        `endif
     `endif
`endif

LUT5    lut_1 (
    .f4    (f[4]),
    .f3    (f[3]),
    .f2    (f[2]),
    .f1    (f[1]),
    .f0    (f[0]),
    .dx    (x1)
`ifdef FM_HACK
    ,.config_data (cfg_data[63:32])
`endif
);
`ifndef CS_FORMALPRO_HACK 
     `ifdef  SIMULATION
//      initial  lut_1.config_data=config_data[63:32];
     `else
        `ifdef FM_HACK
        //BLANK param
        `else
            defparam lut_1.config_data=cfg_data[63:32];
        `endif
     `endif
`endif

assign    x = x1;

MUX2S_L mux_xy (
    .sel    (mode_sel),
    .i0    (x0),
    .i1    (x1),
    .o    (xy) 
);

`ifndef CS_FORMALPRO_HACK 
     `ifdef  SIMULATION
      initial  mux_mode_sel.SEL=mode;
     `else
        `ifdef FM_HACK
        //BLANK param
        `else
            defparam mux_mode_sel.SEL=mode;
        `endif
     `endif
`endif
CFGMUX2S1 mux_mode_sel (
    .i0    (f[5]),
    .i1    (1'b0),
    .o    (mode_sel) 
`ifdef FM_HACK
    ,.SEL (mode)
`endif
);

`endif

endmodule


module FIFOCTRL18KV1(
    rst_n,
    rd_req_n,
    wr_req_n,
	write_drop,
	write_save,
	wrdp_rd_flag,
    clka,
    clkb,
    full,
    empty,
    wptr, 
    rptr,
    wr_mem_n,            
    rd_mem_n,
    overflow,
    underflow,
	prog_full,
	prog_empty,
	peek_en,
	peek_rd_en 
`ifdef FM_HACK
    ,USR_PF
    ,USR_PE
    ,PEEK_MODE
    ,FIFO_EN
    ,R_WIDTH
    ,W_WIDTH
    ,DEPTH_EXT_MODE
`endif
    );


input               rst_n;                  
input               rd_req_n;                
input               wr_req_n;                
input               clka;//read clock
input               clkb;//write clock
input				write_drop;
input				write_save;

output				wrdp_rd_flag;
output              full;
output              empty;
output				prog_full;
output				prog_empty;
output  [13:0] wptr; 
output  [13:0] rptr;
output              wr_mem_n;
output              rd_mem_n;

output              overflow;
output              underflow;//high-active
output				peek_en;
output				peek_rd_en;

`ifdef FM_HACK
    input  [13:0]  USR_PF;
    input  [13:0]  USR_PE;
    input          PEEK_MODE;
    input          FIFO_EN;
    input  [3:0]   R_WIDTH;
    input  [3:0]   W_WIDTH;
    input  [1:0]   DEPTH_EXT_MODE;
`else
    parameter      USR_PF         = 14'b0;
    parameter      USR_PE         = 14'b0;
    parameter      PEEK_MODE      = 1'b0;
    parameter      FIFO_EN        = 1'b0;
    parameter      R_WIDTH        = 4'b0;
    parameter      W_WIDTH        = 4'b0;
    parameter      DEPTH_EXT_MODE = 2'b00;//11 - 18k / 01 - 9k  / others - 4.5k
`endif

`ifndef FM_HACK
    reg gbl_clear_b=1;
    wire GSR;
    glbsr inst( .GSR( GSR )) ;

    initial begin
        gbl_clear_b = 1'b0;
        @(posedge GSR);
        gbl_clear_b = 1'b1;
    end
`else
    wire gbl_clear_b=1;
`endif

/*
   width definition:
   0000=18(16)bit
   1000=9(8)bit
   1100=4bit
   1110=2bit
   1111=1bit
 */

wire			rd_pk,rd_n_m,wr_n_s;
wire			empty_s,empty_m;
wire			underflow_m,overflow_s,underflow_s;
wire			rd_mem_pk,rd_mem_n_m;
//gclk_clk_and clka_gating ( .ck_i0(FIFO_EN), .ck_i1(clka), .ck_out(clka_t));
//gclk_clk_and clkb_gating ( .ck_i0(FIFO_EN), .ck_i1(clkb), .ck_out(clkb_t));

assign clka_t = clka & FIFO_EN;
assign clkb_t = clkb & FIFO_EN;

assign rd_pk = PEEK_MODE ? rd_n_m : rd_req_n;
assign rd_mem_n = PEEK_MODE ? rd_mem_pk : rd_mem_n_m;
assign rd_mem_pk = rd_req_n & rd_mem_n_m;
assign empty = PEEK_MODE ? empty_s : empty_m;
assign underflow = PEEK_MODE ? underflow_s : underflow_m;
// VPERL: GENERATED_BEG

wire rst_n_t = rst_n & gbl_clear_b;

fifo_ctrl_core u_fifo_ctrl_core (
	.w_width	(W_WIDTH[3:0]),
	.r_width	(R_WIDTH[3:0]),
	.depth_ext_mode	(DEPTH_EXT_MODE),
	.peek_mode	(PEEK_MODE),
	.wclk		(clkb_t),
	.rclk		(clka_t),
	.wrst_n		(rst_n_t),
	.rrst_n		(rst_n_t),
	.wr_req_n	(wr_req_n),
	.write_drop	(write_drop),
	.write_save	(write_save),
	.wrdp_rd_flag	(wrdp_rd_flag),
	.rd_req_n	(rd_pk),
	.usr_pf		(USR_PF[13:0]),
	.usr_pe		(USR_PE[13:0]),

	.full		(full),
	.empty		(empty_m),
	.prog_full	(prog_full),
	.prog_empty	(prog_empty),
	.overflow	(overflow),
	.underflow	(underflow_m),
	.wr_mem_n	(wr_mem_n),
	.rd_mem_n	(rd_mem_n_m),
	.wr_addr	(wptr[13:0]),
	.rd_addr	(rptr[13:0]) 
);
// VPERL: GENERATED_END
fifo_pkslice u_fifo_pkslice (
	.clk		(clka_t),
	.rst_n		(rst_n_t),
	.wr_req_n	(wr_n_s),
	.rd_req_n	(rd_req_n),
	.full		(full_s),
	.afull		(afull_s),
	.empty		(empty_s),
	.overflow	(overflow_s),
	.underflow	(underflow_s),
	.wr_en		(peek_en),
	.rd_en		(peek_rd_en)
	);
fifo_pkarbit u_fifo_pkarbit (
	.clk		(clka_t),
	.rst_n		(rst_n_t),
	.empty_m	(empty_m),
	.full_s		(full_s),
	.afull_s	(afull_s),
	.rd_n_m		(rd_n_m),
	.wr_n_s		(wr_n_s),
	.rd_req_usr	(rd_req_n)
	);
endmodule

module hpc_d2s (
	HPC_CLK,
	HPC_CLK_IN,
	HPC_CLK_IP 
`ifdef FM_HACK
	,EN
`endif
);

output		HPC_CLK;
input		HPC_CLK_IN;
input		HPC_CLK_IP;

`ifdef FM_HACK
    input   EN;
`else
    parameter    EN = 1'b0;
`endif

wire		dangling;
assign HPC_CLK  = EN & HPC_CLK_IP;
assign dangling = EN & HPC_CLK_IN;

endmodule

module hpc_s2d (
	HPC_CLK_ON,
	HPC_CLK_OP,
	HPC_CLK 
`ifdef FM_HACK
	,EN
`endif
);

output	HPC_CLK_ON;
output	HPC_CLK_OP;
input	HPC_CLK;

`ifdef FM_HACK
    input  EN;
`else
    parameter    EN = 1'b0;
`endif

assign HPC_CLK_OP  = EN &  HPC_CLK;
assign HPC_CLK_ON  = EN & ~HPC_CLK;

endmodule

module IOC_CMOS(
     clk_en
    ,oen
    ,f_oen
    ,od
    ,f_od
    ,id
    ,f_id
    ,fclk
    ,rstn
    ,setn
`ifdef FM_HACK
    ,CFG_CLK_INV
    ,CFG_DDR
    ,CFG_FOEN_SELN
    ,CFG_FOUT_SELN
    ,CFG_FIN_SELN
    ,CFG_FCLK_GATE_EN
    ,CFG_SETN_INV
    ,CFG_SETN_SYNC
    ,CFG_OEN_SETN_EN
    ,CFG_OD_SETN_EN
    ,CFG_ID_SETN_EN
    ,CFG_RSTN_INV
    ,CFG_RSTN_SYNC
    ,CFG_OEN_RSTN_EN
    ,CFG_OD_RSTN_EN
    ,CFG_ID_RSTN_EN
    ,CFG_DDR_REG
    ,CFG_DDR_PREG
    ,CFG_DDR_NREG
`endif
);

input          clk_en;
input          oen;
output         f_oen;
input  [1:0]   od;
output         f_od;
input          id;
output [1:0]   f_id;
input          fclk;
input          rstn;
input          setn;
`ifdef FM_HACK
input          CFG_CLK_INV;
input          CFG_DDR;
input          CFG_FOEN_SELN;
input          CFG_FOUT_SELN;
input          CFG_FIN_SELN;
input          CFG_FCLK_GATE_EN;
input          CFG_SETN_INV;
input          CFG_SETN_SYNC;
input          CFG_OEN_SETN_EN;
input          CFG_OD_SETN_EN;
input          CFG_ID_SETN_EN;
input          CFG_RSTN_INV;
input          CFG_RSTN_SYNC;
input          CFG_OEN_RSTN_EN;
input          CFG_OD_RSTN_EN;
input          CFG_ID_RSTN_EN;
input          CFG_DDR_REG;
input          CFG_DDR_PREG;
input          CFG_DDR_NREG;
`else
parameter   CFG_CLK_INV                =1'b0;
parameter   CFG_DDR                    =1'b0;
parameter   CFG_FOEN_SELN              =1'b0;
parameter   CFG_FOUT_SELN              =1'b0;
parameter   CFG_FIN_SELN               =1'b0;
parameter   CFG_FCLK_GATE_EN           =1'b0;
parameter   CFG_SETN_INV               =1'b0;
parameter   CFG_SETN_SYNC              =1'b0;
parameter   CFG_OEN_SETN_EN            =1'b0;
parameter   CFG_OD_SETN_EN             =1'b0;
parameter   CFG_ID_SETN_EN             =1'b0;
parameter   CFG_RSTN_INV               =1'b0;
parameter   CFG_RSTN_SYNC              =1'b0;
parameter   CFG_OEN_RSTN_EN            =1'b0;
parameter   CFG_OD_RSTN_EN             =1'b0;
parameter   CFG_ID_RSTN_EN             =1'b0;
parameter   CFG_DDR_REG                =1'b0;
parameter   CFG_DDR_PREG               =1'b0;
parameter   CFG_DDR_NREG               =1'b0;
`endif
`ifndef FM_HACK
    reg cf_rstn;
    wire GSR;
    glbsr inst( .GSR( GSR )) ;

    initial begin
        cf_rstn = 1'b0;
        @(posedge GSR);
        cf_rstn = 1'b1;
    end
`else
    wire cf_rstn = 1'b1;
`endif
wire [1:0] f_id;
wire [1:0] f_id_n;
wire rstn_inv_cfg = CFG_RSTN_INV ? ~rstn : rstn;
wire setn_inv_cfg = CFG_SETN_INV ? ~setn : setn;

//wire fclk_gate_en;
wire fclk_gate_mux;


ioc_latn_ar rstn_syn (
     .ck    (fclk_gate_mux )
    ,.d     (rstn_inv_cfg  )
    ,.q     (rstn_lat      )
    ,.rstn  (cf_rstn       )
);

ioc_latn_ar setn_syn (
     .ck    (fclk_gate_mux )
    ,.d     (setn_inv_cfg  )
    ,.q     (setn_lat      )
    ,.rstn  (cf_rstn       )
);

assign rstn_reg_mux = CFG_RSTN_SYNC ? ~fclk_gate_mux | rstn_lat : rstn_inv_cfg;
assign setn_reg_mux = CFG_SETN_SYNC ? ~fclk_gate_mux | setn_lat : setn_inv_cfg;

assign oen_rstn = CFG_OEN_RSTN_EN ? rstn_reg_mux : 1'b1;
assign od_rstn  = CFG_OD_RSTN_EN ? rstn_reg_mux : 1'b1;
assign id_rstn  = CFG_ID_RSTN_EN ? rstn_reg_mux : 1'b1;

assign t_oen_setn = CFG_OEN_SETN_EN ? setn_reg_mux : 1'b1;
assign t_od_setn  = CFG_OD_SETN_EN ? setn_reg_mux : 1'b1;
assign t_id_setn  = CFG_ID_SETN_EN ? setn_reg_mux : 1'b1;

assign oen_setn = cf_rstn & t_oen_setn;
assign od_setn  = cf_rstn & t_od_setn;
assign id_setn  = cf_rstn & t_id_setn;

assign fclk_cfginv = CFG_CLK_INV ? ~fclk : fclk;
//clk_inv u_fclk_inv ( .ck_(fclk), .ck_n(fclk_inv));
//gclk_clk_mux u_fclk_cfginv (.ck_i0(fclk), .ck_i1(fclk_inv), .sel(CFG_CLK_INV), .ck_out(fclk_cfginv));

reg fclk_gate_en;
always@(*)
begin
    if (CFG_FCLK_GATE_EN)
        fclk_gate_en <= 1'b1;
    else
    begin
        if (!fclk_cfginv)
            fclk_gate_en <= clk_en;
        else
            fclk_gate_en <= fclk_gate_en;
    end
end
assign fclk_gate_mux = fclk_gate_en & fclk_cfginv;

//assign CFG_FCLK_GATE_EN_inv = ~CFG_FCLK_GATE_EN;
//LNSNQD4BWP u0_fclk_gate (.EN(fclk_cfginv),.D(clk_en),.SDN(CFG_FCLK_GATE_EN_inv),.Q(fclk_gate_en));
//gclk_clk_and u_fclk_gate (.ck_i0(fclk_cfginv),.ck_i1(fclk_gate_en),.ck_out(fclk_gate_mux));

//ECO 20140521 beg
//assign ioc_clk_out = fclk_gate_mux;
//ECO 20140521 end

//f_oen
ioc_dff_asr u0_oen(
     .ck     ( fclk_gate_mux )
    ,.d      ( oen           )
    ,.q      ( oen_reg       )
    ,.rstn   ( oen_rstn      )
    ,.setn   ( oen_setn      )
);

assign f_oen = (CFG_FOEN_SELN == 0) ? oen_reg : oen;

//f_od
ioc_dff_asr u_od0(
     .ck     ( fclk_gate_mux )
    ,.d      ( od[0]        )
    ,.q      ( out_reg0      )
    ,.rstn   ( od_rstn       )
    ,.setn   ( od_setn       )
);

ioc_dff_asr u_od1(
     .ck     ( fclk_gate_mux )
    ,.d      ( od[1]        )
    ,.q      ( out_reg1      )
    ,.rstn   ( od_rstn       )
    ,.setn   ( od_setn       )
);
assign oddr_reg0 = CFG_DDR_REG ? out_reg0 : od[0];
assign oddr_reg1 = CFG_DDR_REG ? out_reg1 : od[1];

ioc_dff_asr u_od2(
     .ck     ( fclk_gate_mux )
    ,.d      ( oddr_reg0     )
    ,.q      ( out_reg2      )
    ,.rstn   ( od_rstn       )
    ,.setn   ( od_setn       )
);

ioc_dffn_asr u_od3(
     .ckb    ( fclk_gate_mux )
    ,.d      ( oddr_reg1     )
    ,.q      ( out_reg3      )
    ,.rstn   ( od_rstn       )
    ,.setn   ( od_setn       )
);
//assign ddr_sel = ~(fclk_gate_mux & CFG_DDR);
assign ddr_sel = fclk_gate_mux & CFG_DDR;
assign f_od_ddr = ddr_sel ? out_reg3 : out_reg2;
assign f_od = (CFG_FOUT_SELN == 0) ? f_od_ddr : od[0];
//assign f_od_fb = f_od;

//f_id
ioc_dff_asr u_id0(
     .ck     ( fclk_gate_mux )
    ,.d      ( id            )
    ,.q      ( iddr_reg0       )
    ,.rstn   ( id_rstn       )
    ,.setn   ( id_setn       )
);

ioc_dffn_asr u_id1(
     .ckb    ( fclk_gate_mux )
    ,.d      ( id            )
    ,.q      ( iddr_reg1       )
    ,.rstn   ( id_rstn       )
    ,.setn   ( id_setn       )
);

ioc_dff_asr u_id2(
     .ck     ( fclk_gate_mux )
    ,.d      ( iddr_reg0     )
    ,.q      ( in_reg0       )
    ,.rstn   ( id_rstn       )
    ,.setn   ( id_setn       )
);

ioc_dff_asr u_id3(
     .ck     ( fclk_gate_mux )
    ,.d      ( iddr_reg1     )
    ,.q      ( in_reg1       )
    ,.rstn   ( id_rstn       )
    ,.setn   ( id_setn       )
);

assign f_id0_t = CFG_DDR_PREG ? in_reg0 : iddr_reg0;
assign f_id[0] = (CFG_FIN_SELN == 0) ? f_id0_t : id;
assign f_id[1] = CFG_DDR_NREG ? in_reg1 : iddr_reg1;

endmodule

module IOC_LVDS (
	//port
	geclk0_up_il,
	geclk0_up_ol,
	rxd_dr,
	txd_out,
	ted_out,
	shiftout0_il,
	shiftout0_ol,
	shiftout1_il,
	shiftout1_ol,
	q,

	oen,
	rxd_in,
	shiftin0_il,
	shiftin0_ol,
	shiftin1_il,
	shiftin1_ol,
	update_il,
	update_b_il,
	update_ol,
	update_b_ol,
	clken,
	rstn,
	setn,
	feclk,
	sclk,
	test,
	d
	//PARAMETER
	`ifdef FM_HACK
	,CFG_CK_INV
	,CFG_CK_PAD_EN
	,CFG_DDR_IN_NREG
	,CFG_DDR_IN_NREG_DFF
	,CFG_DDR_IN_PREG
	,CFG_DDR_IN_PREG_DFF
	,CFG_DDR_OUT
	,CFG_DDR_OUT_REG
	,CFG_DQS_CLK
	,CFG_ECLK_INV
	,CFG_FASTIN
	,CFG_FCLK0_I_EN
	,CFG_FCLK0_OEN
	,CFG_FCLK0_O_EN
	,CFG_FCLK0_RS_EN
	,CFG_FCLK0_UPI_EN
	,CFG_FCLK0_UPO_EN
	,CFG_FCLK1_I_EN
	,CFG_FCLK1_O_EN
	,CFG_FCLK_INV
	,CFG_FOUT_SEL
	,CFG_GEAR_IN
	,CFG_GEAR_OUT
	,CFG_GECLK0_I_EN
	,CFG_GECLK0_O_EN
	,CFG_GECLK1_I_EN
	,CFG_GECLK1_O_EN
	,CFG_GSCLK0_I_EN
	,CFG_GSCLK0_O_EN
	,CFG_GSCLK1_I_EN
	,CFG_GSCLK1_O_EN
	,CFG_IN_EN
	,CFG_OEN_INV
	,CFG_OEN_SEL
	,CFG_OFDBK
	,CFG_OUT_SEL
	,CFG_RSTN
	,CFG_SCLK_INV
	,CFG_SETN
	,CFG_SLAVE_IN
	,CFG_TEST
	`endif
	);
output	geclk0_up_il;
output	geclk0_up_ol;
output	rxd_dr;
output	txd_out;
output	ted_out;
output	shiftout0_il;
output	shiftout0_ol;
output	shiftout1_il;
output	shiftout1_ol;
output	[7:0]	q;

input	oen;
input	rxd_in;
input	shiftin0_il;
input	shiftin0_ol;
input	shiftin1_il;
input	shiftin1_ol;
input	update_il;
input	update_b_il;
input	update_ol;
input	update_b_ol;
input	clken;
input	rstn;
input	setn;
input	feclk;
input	sclk;
input	[7:0]	test;
input	[7:0]	d;
`ifdef FM_HACK
input	CFG_CK_INV;
input	CFG_CK_PAD_EN;
input	CFG_DDR_IN_NREG;
input	CFG_DDR_IN_NREG_DFF;
input	CFG_DDR_IN_PREG;
input	CFG_DDR_IN_PREG_DFF;
input	CFG_DDR_OUT;
input	CFG_DDR_OUT_REG;
input	CFG_DQS_CLK;
input	CFG_ECLK_INV;
input	CFG_FASTIN;
input	CFG_FCLK0_I_EN;
input	CFG_FCLK0_OEN;
input	CFG_FCLK0_O_EN;
input	CFG_FCLK0_RS_EN;
input	CFG_FCLK0_UPI_EN;
input	CFG_FCLK0_UPO_EN;
input	CFG_FCLK1_I_EN;
input	CFG_FCLK1_O_EN;
input	CFG_FCLK_INV;
input	CFG_FOUT_SEL;
input	CFG_GEAR_OUT;
input	CFG_GECLK0_I_EN;
input	CFG_GECLK0_O_EN;
input	CFG_GECLK1_I_EN;
input	CFG_GECLK1_O_EN;
input	CFG_GSCLK0_I_EN;
input	CFG_GSCLK0_O_EN;
input	CFG_GSCLK1_I_EN;
input	CFG_GSCLK1_O_EN;
input	CFG_OEN_INV;
input	CFG_OFDBK;
input	CFG_SCLK_INV;
input	CFG_SLAVE_IN;
input	[7:0]	CFG_GEAR_IN;
input	[1:0]	CFG_IN_EN;
input	[3:0]	CFG_OEN_SEL;
input	[2:0]	CFG_OUT_SEL;
input	[4:0]	CFG_RSTN;
input	[4:0]	CFG_SETN;
input	[7:0]	CFG_TEST;
`else
parameter	CFG_CK_INV=1'b0;
parameter	CFG_CK_PAD_EN=1'b0;
parameter	CFG_DDR_IN_NREG=1'b0;
parameter	CFG_DDR_IN_NREG_DFF=1'b0;
parameter	CFG_DDR_IN_PREG=1'b0;
parameter	CFG_DDR_IN_PREG_DFF=1'b0;
parameter	CFG_DDR_OUT=1'b0;
parameter	CFG_DDR_OUT_REG=1'b0;
parameter	CFG_DQS_CLK=1'b0;
parameter	CFG_ECLK_INV=1'b0;
parameter	CFG_FASTIN=1'b0;
parameter	CFG_FCLK0_I_EN=1'b0;
parameter	CFG_FCLK0_OEN=1'b0;
parameter	CFG_FCLK0_O_EN=1'b0;
parameter	CFG_FCLK0_RS_EN=1'b0;
parameter	CFG_FCLK0_UPI_EN=1'b0;
parameter	CFG_FCLK0_UPO_EN=1'b0;
parameter	CFG_FCLK1_I_EN=1'b0;
parameter	CFG_FCLK1_O_EN=1'b0;
parameter	CFG_FCLK_INV=1'b0;
parameter	CFG_FOUT_SEL=1'b0;
parameter	CFG_GEAR_OUT=1'b0;
parameter	CFG_GECLK0_I_EN=1'b0;
parameter	CFG_GECLK0_O_EN=1'b0;
parameter	CFG_GECLK1_I_EN=1'b0;
parameter	CFG_GECLK1_O_EN=1'b0;
parameter	CFG_GSCLK0_I_EN=1'b0;
parameter	CFG_GSCLK0_O_EN=1'b0;
parameter	CFG_GSCLK1_I_EN=1'b0;
parameter	CFG_GSCLK1_O_EN=1'b0;
parameter	CFG_OEN_INV=1'b0;
parameter	CFG_OFDBK=1'b0;
parameter	CFG_SCLK_INV=1'b0;
parameter	CFG_SLAVE_IN=1'b0;
parameter	CFG_GEAR_IN=8'b0;
parameter	CFG_IN_EN=2'b0;
parameter	CFG_OEN_SEL=4'b0;
parameter	CFG_OUT_SEL=3'b0;
parameter	CFG_RSTN=5'b0;
parameter	CFG_SETN=5'b0;
parameter	CFG_TEST=8'b0;
`endif
wire	[7:0]	CFG_GEAR_IN_              = ~CFG_GEAR_IN;
wire	[1:0]	CFG_IN_EN_                = ~CFG_IN_EN;
wire	[2:0]	CFG_OUT_SEL_              = ~CFG_OUT_SEL;
wire	[4:0]	CFG_RSTN_                 = ~CFG_RSTN;
wire	[4:0]	CFG_SETN_                 = ~CFG_SETN;
wire	[7:0]	CFG_TEST_                 = ~CFG_TEST;
wire			CFG_CK_INV_               = ~CFG_CK_INV;
wire			CFG_DDR_IN_NREG_          = ~CFG_DDR_IN_NREG;
wire			CFG_DDR_IN_NREG_DFF_      = ~CFG_DDR_IN_NREG_DFF;
wire			CFG_DDR_IN_PREG_          = ~CFG_DDR_IN_PREG;
wire			CFG_DDR_IN_PREG_DFF_      = ~CFG_DDR_IN_PREG_DFF;
wire			CFG_DDR_OUT_REG_          = ~CFG_DDR_OUT_REG;
wire			CFG_DQS_CLK_              = ~CFG_DQS_CLK;
wire			CFG_FASTIN_               = ~CFG_FASTIN;
wire			CFG_FOUT_SEL_             = ~CFG_FOUT_SEL;
wire			CFG_GEAR_OUT_             = ~CFG_GEAR_OUT;
wire			CFG_OEN_INV_              = ~CFG_OEN_INV;
wire			CFG_OFDBK_                = ~CFG_OFDBK;
wire			CFG_SLAVE_IN_             = ~CFG_SLAVE_IN;
`ifndef FM_HACK
reg gbl_clear_b;
wire GSR;
glbsr inst( .GSR( GSR )) ;

initial begin
gbl_clear_b = 1'b0;
@(posedge GSR);
gbl_clear_b = 1'b1;
end
`else
wire gbl_clear_b = 1'b1;
`endif

assign rxd_dr = CFG_CK_PAD_EN & rxd_in;
wire	txd_in,txd_in_b;
assign txd_in_b = ~txd_in;
assign txd_out =	({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b001_110) ? 1'b0 :
					({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b010_101) ? txd_in_b :
					({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b100_011) ? txd_in :
					({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b000_111) ? 1'b1 : 1'bx;
wire	datain;
assign datain =	({CFG_OFDBK,CFG_OFDBK_} == 2'b01) ? rxd_in :
				({CFG_OFDBK,CFG_OFDBK_} == 2'b10) ? txd_in : 1'bx;
// VPERL: GENERATED_BEG


CLK Iclk (
	.CFG_CKEN_INV		(CFG_CK_INV),
	.CFG_CKEN_INV_		(CFG_CK_INV_),
	.CFG_FCLK0_I_EN		(CFG_FCLK0_I_EN),
	.CFG_FCLK0_OEN		(CFG_FCLK0_OEN),
	.CFG_FCLK0_O_EN		(CFG_FCLK0_O_EN),
	.CFG_FCLK0_RS_EN	(CFG_FCLK0_RS_EN),
	.CFG_FCLK0_UPI_EN	(CFG_FCLK0_UPI_EN),
	.CFG_FCLK0_UPO_EN	(CFG_FCLK0_UPO_EN),
	.CFG_FCLK1_I_EN		(CFG_FCLK1_I_EN),
	.CFG_FCLK1_O_EN		(CFG_FCLK1_O_EN),
	.CFG_GECLK0_I_EN	(CFG_GECLK0_I_EN),
	.CFG_GECLK0_O_EN	(CFG_GECLK0_O_EN),
	.CFG_GECLK1_I_EN	(CFG_GECLK1_I_EN),
	.CFG_GECLK1_O_EN	(CFG_GECLK1_O_EN),
	.CFG_GSCLK0_I_EN	(CFG_GSCLK0_I_EN),
	.CFG_GSCLK0_O_EN	(CFG_GSCLK0_O_EN),
	.CFG_GSCLK1_I_EN	(CFG_GSCLK1_I_EN),
	.CFG_GSCLK1_O_EN	(CFG_GSCLK1_O_EN),
	.CFG_RSTN_ID_EN		(CFG_RSTN[4]),
	.CFG_RSTN_ID_EN_	(CFG_RSTN_[4]),
	.CFG_RSTN_INV		(CFG_RSTN[1]),
	.CFG_RSTN_INV_		(CFG_RSTN_[1]),
	.CFG_RSTN_OD_EN		(CFG_RSTN[3]),
	.CFG_RSTN_OD_EN_	(CFG_RSTN_[3]),
	.CFG_RSTN_OEN_EN	(CFG_RSTN[2]),
	.CFG_RSTN_OEN_EN_	(CFG_RSTN_[2]),
	.CFG_RSTN_SYNC		(CFG_RSTN[0]),
	.CFG_RSTN_SYNC_		(CFG_RSTN_[0]),
	.CFG_SETN_ID_EN		(CFG_SETN[4]),
	.CFG_SETN_ID_EN_	(CFG_SETN_[4]),
	.CFG_SETN_INV		(CFG_SETN[1]),
	.CFG_SETN_INV_		(CFG_SETN_[1]),
	.CFG_SETN_OD_EN		(CFG_SETN[3]),
	.CFG_SETN_OD_EN_	(CFG_SETN_[3]),
	.CFG_SETN_OEN_EN	(CFG_SETN[2]),
	.CFG_SETN_OEN_EN_	(CFG_SETN_[2]),
	.CFG_SETN_SYNC		(CFG_SETN[0]),
	.CFG_SETN_SYNC_		(CFG_SETN_[0]),
	.CFG_SCLK_INV		(CFG_SCLK_INV),
	.CFG_ECLK_INV		(CFG_ECLK_INV),
	.setn			(setn),
	.rstn			(rstn),
	.clk_en			(clken),
	.sclk			(sclk),
	.feclk			(feclk),

	.fclk0_il		(fclk0_il),
	.fclk0_oen		(oen_fclk0),
	.fclk0_ol		(fclk0_ol),
	.fclk1_il		(fclk1_il),
	.fclk1_ol		(fclk1_ol),
	.geclk0_il		(geclk0_il),
	.geclk0_ol		(geclk0_ol),
	.geclk0_up_il		(geclk0_up_il),
	.geclk0_up_ol		(geclk0_up_ol),
	.geclk1_il		(geclk1_il),
	.geclk1_ol		(geclk1_ol),
	.gsclk0_il		(gsclk0_il),
	.gsclk0_ol		(gsclk0_ol),
	.gsclk1_il		(gsclk1_il),
	.gsclk1_ol		(gsclk1_ol),
	.id_rst			(id_rst),
	.id_setn		(id_set_),
	.od_rst			(od_rst),
	.od_setn		(od_set_),
	.oen_rst		(oen_rst),
	.oen_setn		(oen_set_) 
);

ILOGIC Iilg (
	.datain			(datain),
	.fclk0			(fclk0_il),
	.fclk1			(fclk1_il),
	.geclk0			(geclk0_il),
	.geclk1			(geclk1_il),
	.gsclk0			(gsclk0_il),
	.gsclk1			(gsclk1_il),
	.init_b			(1'b1),
	.rst			(id_rst),
	.set_			(id_set_),
	.shiftin0		(shiftin0_il),
	.shiftin1		(shiftin1_il),
	.update			(update_il),
	.update_		(update_b_il),
	.usermode		(gbl_clear_b),
	.test			(test[7:0]),
	.CFG_DDR_IN_NREG	(CFG_DDR_IN_NREG),
	.CFG_DDR_IN_NREG_DFF	(CFG_DDR_IN_NREG_DFF),
	.CFG_DDR_IN_PREG	(CFG_DDR_IN_PREG),
	.CFG_DDR_IN_PREG_DFF	(CFG_DDR_IN_PREG_DFF),
	.CFG_DQS_CLK		(CFG_DQS_CLK),
	.CFG_FASTIN		(CFG_FASTIN),
	.CFG_SLAVE_IN		(CFG_SLAVE_IN),
	.CFG_TEST		(CFG_TEST[7:0]),
	.CFG_IN_EN		(CFG_IN_EN[1:0]),
	.CFG_GEAR_IN		(CFG_GEAR_IN[7:0]),
	.CFG_DDR_IN_NREG_	(CFG_DDR_IN_NREG_),
	.CFG_DDR_IN_NREG_DFF_	(CFG_DDR_IN_NREG_DFF_),
	.CFG_DDR_IN_PREG_	(CFG_DDR_IN_PREG_),
	.CFG_DDR_IN_PREG_DFF_	(CFG_DDR_IN_PREG_DFF_),
	.CFG_DQS_CLK_		(CFG_DQS_CLK_),
	.CFG_FASTIN_		(CFG_FASTIN_),
	.CFG_SLAVE_IN_		(CFG_SLAVE_IN_),
	.CFG_TEST_		(CFG_TEST_[7:0]),
	.CFG_IN_EN_		(CFG_IN_EN_[1:0]),
	.CFG_GEAR_IN_		(CFG_GEAR_IN_[7:0]),

	.shiftout0		(shiftout0_il),
	.shiftout1		(shiftout1_il),
	.dataout		(q[7:0]) 
);

OLOGIC Iolg (
	.fclk0			(fclk0_ol),
	.fclk1			(fclk1_ol),
	.geclk0			(geclk0_ol),
	.geclk1			(geclk1_ol),
	.gsclk0			(gsclk0_ol),
	.gsclk1			(gsclk1_ol),
	.rst			(od_rst),
	.set_			(od_set_),
	.shiftin0		(shiftin0_ol),
	.shiftin1		(shiftin1_ol),
	.update			(update_ol),
	.update_		(update_b_ol),
	.usermode		(gbl_clear_b),
	.datain			(d[7:0]),
	.CFG_DDR_OUT		(CFG_DDR_OUT),
	.CFG_DDR_OUT_REG	(CFG_DDR_OUT_REG),
	.CFG_DDR_OUT_REG_	(CFG_DDR_OUT_REG_),
	.CFG_FCLK_INV		(CFG_FCLK_INV),
	.CFG_FOUT_SEL		(CFG_FOUT_SEL),
	.CFG_FOUT_SEL_		(CFG_FOUT_SEL_),
	.CFG_GEAR_OUT		(CFG_GEAR_OUT),
	.CFG_GEAR_OUT_		(CFG_GEAR_OUT_),

	.dataout		(txd_in),
	.shiftout0		(shiftout0_ol),
	.shiftout1		(shiftout1_ol) 
);

OENC Ioen (
	.clk		(oen_fclk0),
	.gbl_clear_b	(gbl_clear_b),
	.init_b		(1'b1),
	.oen		(oen),
	.rst		(oen_rst),
	.set_		(oen_set_),
	.CFG_OEN_INV	(CFG_OEN_INV),
	.CFG_OEN_INV_	(CFG_OEN_INV_),
	.CFG_OEN_SEL	(CFG_OEN_SEL[3:0]),

	.f_oen		(ted_out) 
);
// VPERL: GENERATED_END
endmodule

module JTAG_DBWV1(
    // Outputs
	jtag_fp_drck     , 
	jtag_fp_reset ,
	jtag_fp_sel,
	jtag_fp_capture,
	jtag_fp_shift,
	jtag_fp_update,
	jtag_fp_tdi      ,
    // Inputs
//	jtag_fp_usermode,
	jtag_fp_tdo
);

    // Outputs
	output jtag_fp_drck     ; 
	output jtag_fp_reset ;
	output [1:0] jtag_fp_sel;
	output jtag_fp_capture;
	output jtag_fp_shift;
	output jtag_fp_update;
	output jtag_fp_tdi      ;
    // Inputs
//	input  jtag_fp_usermode;
	input  jtag_fp_tdo;
    
endmodule
//----------------------------------------------------------------------------
//
// module: LBUF
//
// description: register control for 8 REGs in LE.
// config:      1 bit enable control
//              1 bit invert sense of "en" input
//              1 bit invert clk control
//              1 bit close clk control
//              1 bit REG or LATCH selection
//              1 bit SYNC or ASYNC set/reset selection
//              1 bit ASYNC set/reset assert even if SYNC is configured (deassert with be synchronized)
//              1 bit ALLOW_SR to enable set/reset (if =0, ignores "sr" input)
//              1 bit invert sense of "sr" input
//
// notes: RST and SET inputs are active high.
//
//----------------------------------------------------------------------------
module LBUF (
        asr,
        mclkb,
        sclk,

        clk,
        en,
        sr
`ifdef FM_HACK
		,CFG_EN       
		,CFG_INV      
		,CFG_HASCLK   
		,CFG_LAT      
		,CFG_SYNC     
		,CFG_ALLOW_SR 
		,CFG_INV_EN   
		,CFG_INV_SR   
`endif
);

output  asr;
output  mclkb;
output  sclk;

input   clk;
input   en;
input   sr;


`ifdef CS_FORMALPRO_HACK
   wire        CFG_EN      ;    // enable clock gating
   wire        CFG_INV     ;    // invert clock input (emulate negedge FFs, using posedge FFs)
   wire        CFG_HASCLK   ;    // allow clock
   wire        CFG_LAT     ;    // if =1, hold master clock "open"
   wire        CFG_SYNC    ;    // synchronize set/reset assert/deassert with active clock
   wire        CFG_ALLOW_SR ;    // allow set/reset; if =0, ignore "sr" input
   wire        CFG_INV_EN ;    // treat "en" input as active-low
   wire        CFG_INV_SR ;    // treat "sr" input as active-low
`else
     `ifdef  SIMULATION
          reg        CFG_EN       = 1'b0;
          reg        CFG_INV      = 1'b0;
          reg        CFG_HASCLK   = 1'b0;
          reg        CFG_LAT      = 1'b0;
          reg        CFG_SYNC     = 1'b0;
          reg        CFG_ALLOW_SR = 1'b0;
          reg        CFG_INV_EN   = 1'b0;
          reg        CFG_INV_SR   = 1'b0;
     `else
		`ifdef FM_HACK
			input  CFG_EN       ;
			input  CFG_INV      ;
			input  CFG_HASCLK   ;
			input  CFG_LAT      ;
			input  CFG_SYNC     ;
			input  CFG_ALLOW_SR ;
			input  CFG_INV_EN   ;
			input  CFG_INV_SR   ;
		`else
			parameter  CFG_EN       = 1'b0;
          	parameter  CFG_INV      = 1'b0;
          	parameter  CFG_HASCLK   = 1'b0;
          	parameter  CFG_LAT      = 1'b0;
          	parameter  CFG_SYNC     = 1'b0;
          	parameter  CFG_ALLOW_SR = 1'b0;
          	parameter  CFG_INV_EN   = 1'b0;
          	parameter  CFG_INV_SR   = 1'b0;
		`endif
     `endif
`endif

reg         en_latch_b;
wire        en_latch;
wire        clk1;
wire        clk2;
wire        sr_ff;

wire GSR;
glbsr inst( .GSR( GSR )) ;

initial begin
    en_latch_b = 1'b0;
    @(posedge GSR);
    en_latch_b = 1'b1;
end

`ifndef CS_SW_SKEL
    assign    clk1 = (CFG_HASCLK == 1'b1)  ?  clk : 1'b1;
    assign    clk2 = (CFG_INV   == 1'b1)  ? !clk1: clk1;

    wire    clkb = ~clk2;

    wire    sri = (CFG_INV_SR == 1'b1) ? ~sr : sr ;
    wire    eni = (CFG_INV_EN == 1'b1) ? ~en : en ;

    wire    allow_sr    = CFG_ALLOW_SR ;    // actually CFG_ALLOW_SR & gbl_cfg_done & gbl_clear_b
    wire    sr_allowed    = allow_sr? sri: 1'b1 ;
    wire    sr_allowed_i  = ~sr_allowed ;
   
    reg sr_latch;

    always @(*) begin
      if (allow_sr == 0) sr_latch <= sr_allowed_i ;	 
      else if (clkb == 1) sr_latch <= sr_allowed_i ;
    end
    
    wire    sync_sr = sr_latch & clk2;

    assign  asr = (CFG_SYNC == 1'b1) ? !sync_sr : sr_allowed ;

    assign  mclkb = (CFG_LAT == 1'b1)? 1'b0 :
                                       (clk2 & en_latch);

    always @(clkb or eni or CFG_EN) begin
       if (clkb == 1) en_latch_b <= !eni;
    end
    assign en_latch = !en_latch_b | ~CFG_EN;

    assign sclk = clk2 & en_latch;


    specify

        ( clk =>  sclk ) = (0,0);


    endspecify


`endif

endmodule

//----------------------------------------------------------------------------
//
// module: LRAM64
//
//----------------------------------------------------------------------------
module LRAM64 (
    x,
    xy,
    shiftout,
    
    di0,
    f,
    we,
    preda,
    predb
`ifdef FM_HACK
    ,mode
    ,config_data
`endif
);

    output x;
    output xy;
    output shiftout;

    input di0;
    input [5:0] f;
    input we;
    input [4:0] preda;
    input [7:0] predb;
    
    `ifdef  SIMULATION
        reg [63:0] config_data = 64'h0000_0000_0000_0000;
        reg [2:0]  mode = 3'b000;
    `else
        `ifdef FM_HACK
            input    [2:0]    mode;
            input    [63:0]    config_data;
        `else
            parameter mode = 3'b000;
            parameter  [63:0] config_data = 64'h0000_0000_0000_0000;
        `endif
    `endif

    initial begin
    # 1;
    if (mode == 3'b110 || mode == 3'b111) begin
        $display("Attribute Syntax Error : The attribute int_mode on LRAM64 instance %m is set to %d.  Legal values for this attribute are 3'b000, 3'b001, 3'b010, 3'b011, 3'b100 or 3'b101.", mode);
        $finish;
    end
    end
    
    `ifdef SIMULATION    
        reg [63:0] cfg_data;
        initial #1 cfg_data = ~config_data;
    `else 
        `ifndef FM_HACK
            localparam [63:0] cfg_data = ~config_data;
        `else
            wire [63:0] cfg_data = ~config_data;
        `endif
    `endif    
    //Begin of FG6X2 logic
    LUT5    lut_0 (
        .f4    (f[4]),
        .f3    (f[3]),
        .f2    (f[2]),
        .f1    (f[1]),
        .f0    (f[0]),
        .dx    (x0)
    `ifdef FM_HACK
        ,.config_data (cfg_data[31:0])
    `endif
    );
    `ifndef CS_FORMALPRO_HACK 
         `ifdef  SIMULATION
          initial  lut_0.config_data=cfg_data[31:0];
         `else
            `ifdef FM_HACK
                
            `else
                defparam lut_0.config_data=cfg_data[31:0];
            `endif
         `endif
    `endif

    LUT5    lut_1 (
        .f4    (f[4]),
        .f3    (f[3]),
        .f2    (f[2]),
        .f1    (f[1]),
        .f0    (f[0]),
        .dx    (x1)
    `ifdef FM_HACK
        ,.config_data (cfg_data[63:32])
    `endif
    );
    `ifndef CS_FORMALPRO_HACK 
         `ifdef  SIMULATION
          initial  lut_1.config_data=cfg_data[63:32];
         `else
            `ifdef FM_HACK

            `else
                defparam lut_1.config_data=cfg_data[63:32];
            `endif
         `endif
    `endif

    assign    fg_6x2_x = x1; 

    wire mux_mode_sel = (mode == 3'b000) ? f[5] : 
                        (mode == 3'b001) ? 1'b0 :
                        mux_mode_sel; 
    
    assign fg_6x2_xy = (mux_mode_sel == 1'b0) ? x0 : 
                       (mux_mode_sel == 1'b1) ? x1 :
                       (x0  == x1  ) ? x0 : 1'bx;
    //End of FG6X2 logic function

    //Begin of LRAM logic function
    wire [31:0] wl;
    wire [31:0] mux_marin_0, mux_marin_1;
    wire [4:0] rdaddr;
    wire lram_x, lram_xy;
    
    reg di0_q;
    reg di1_q;
    
    reg [1:0] mar [31:0];
    
    reg lram_doutx;
    reg lram_doutxy;
    
    integer lram_count;
    
    initial begin
    #1;
    for(lram_count = 0; lram_count <32; lram_count = lram_count + 1) begin
            mar[lram_count] = {cfg_data[lram_count + 32], cfg_data[lram_count]};
        end
    end
    
    //word line decoder
    genvar i;
    generate
        for(i = 0; i < 32; i = i + 1) begin: wl_decoder
            assign wl[i] = preda[i%4] && predb[i/4] && we;
        end
    endgenerate
    
    //f[5] input select
    wire muxf5_o0 = (mode == 3'b010) ? f[5] : 
                    (mode == 3'b011) ? muxf5_o0 :
                    muxf5_o0;
    wire muxf5_o1 = (mode == 3'b011) ? f[5] : 
                    (mode == 3'b010) ? muxf5_o1 :
                    muxf5_o1;
    
    //data input registers
    always @ (posedge we) begin
        di0_q <= di0;
        di1_q <= muxf5_o1;
    end
    
    wire wr_muxsel = (mode == 3'b010) ? preda[4] :
                     (mode == 3'b011) ? 1'b0 :
                     wr_muxsel;
    wire muxdi0_o0 = (wr_muxsel == 0) ? di0_q : muxdi0_o0;
    wire muxdi0_o1 = (wr_muxsel == 1) ? di0_q : muxdi0_o1;
    
    wire muxdi1_o = (mode == 3'b011) ? di1_q : 
                    (mode == 3'b010) ? muxdi0_o1 :
                    muxdi1_o;

    //MAR input MUXs
    genvar j;
    generate
        for(j = 0; j < 32; j = j + 1) begin: marin_mux
            assign mux_marin_0[j] = (mode == 3'b011) ? muxdi0_o0 :
                    (preda[4] == 0) ? muxdi0_o0 : 
                    mar[j][0];
            assign mux_marin_1[j] = (mode == 3'b011) ? muxdi1_o :
                    (preda[4] == 1) ? muxdi1_o : 
                    mar[j][1];
        end
    endgenerate
    
    //MAR latches
    genvar k;
    generate
    for(k = 0; k < 32; k = k + 1) begin: mar_latches
        always @ (mux_marin_1[k] or mux_marin_0[k] or wl[k]) begin
            if (wl[k] == 1'b1)
                 mar[k] <= {mux_marin_1[k], mux_marin_0[k]};
        end    
    end
    endgenerate
    
    wire lram_muxsel = (mode == 3'b011) ? 1'b0 : 
                       (mode == 3'b010) ? muxf5_o0 :
                       lram_muxsel;
    
    assign rdaddr = f[4:0]; 

    always @ (*) begin
        {lram_doutx, lram_doutxy} = mar[rdaddr];
    end
    wire lram_muxxy = (lram_muxsel == 1'b0) ? lram_doutxy : 
                      (lram_muxsel == 1'b1) ? lram_doutx :
                      1'bx;
    
    assign lram_x = lram_doutx;
    assign lram_xy = lram_muxxy;
    
    //End of LRAM logic function
    
    
    //Begin of SR logic function
    reg [15:0] dataxy, datax;
    reg sr_doutx, sr_doutxy;
    
    wire shiftin0, shiftin1;
    wire [3:0] raddr;
    
    integer sr_count, sr_baseaddrr;    
    initial begin
    # 1;
        for(sr_count = 0; sr_count <16; sr_count = sr_count + 1) begin
            sr_baseaddrr = sr_count * 2 + 1;
            dataxy[sr_count] = cfg_data[sr_baseaddrr];
            datax[sr_count] = cfg_data[sr_baseaddrr + 32];
        end
    end    
    
    wire mux_shift1 = (mode == 3'b101) ? f[5] : 
                      (mode == 3'b100) ? dataxy[15] :
                      mux_shift1;
    assign shiftin0 = di0;
    assign shiftin1 = mux_shift1;
    
    always @(posedge we) begin
        {dataxy[15:0]} <= {dataxy[14:0], shiftin0};
        {datax[15:0]} <= {datax[14:0], shiftin1};
    end
    
    assign raddr = f[4:1];
    always @ (*) begin
        {sr_doutx, sr_doutxy} = {datax[raddr], dataxy[raddr]};
    end
    
    wire sr_muxsel = (mode == 3'b101) ? 1'b0 : 
                     (mode == 3'b100) ? f[5] :
                     sr_muxsel;
    wire sr_muxxy = (sr_muxsel == 1'b0) ? sr_doutxy : 
                    (sr_muxsel == 1'b1) ? sr_doutx :
                    1'bx;

    assign sr_x = sr_doutx;
    assign sr_xy = sr_muxxy;
    
    assign x = (mode == 3'b000) ? fg_6x2_x :
               (mode == 3'b001) ? fg_6x2_x :
               (mode == 3'b011) ? lram_x :
               (mode == 3'b010) ? lram_x :
               (mode == 3'b100) ? sr_x :
               (mode == 3'b101) ? sr_x :
               1'bx;
    assign xy = (mode == 3'b000) ? fg_6x2_xy :
                (mode == 3'b001) ? fg_6x2_xy :
                (mode == 3'b011) ? lram_xy :
                (mode == 3'b010) ? lram_xy :
                (mode == 3'b100) ? sr_xy :
                (mode == 3'b101) ? sr_xy :
                1'bx;
    
    assign shiftout = datax[15];

endmodule

//----------------------------------------------------------------------------
//
// module: LRAM_CTRL
//
//----------------------------------------------------------------------------
module LRAM_CTRL (
    weq0,        //output gated clocks to each LRAM64
    weq1,
    weq2,
    weq3,
    preda,        //pre-decoder outputs to all 4 LRAM64s
    predb,
    
    clk0,        //input gated clocks from PLBBUF
    clk1,
    wa            //input write address from xbar
`ifdef FM_HACK
	,we_mode
	,clksel
`endif
);

    output weq0;
    output weq1;
    output weq2;
    output weq3;
    output [4:0] preda;        //preda[4] = wa[5]
    output [7:0] predb;

    input clk0;
    input clk1;
    input [7:0] wa;
	
    `ifdef  SIMULATION
		reg [1:0] we_mode = 2'b00;
		reg [1:0] clksel = 2'b00;
    `else
		`ifdef FM_HACK
			input	[1:0]	we_mode;
			input	[1:0]	clksel;
		`else
	        	parameter we_mode = 2'b00;
		        parameter clksel = 2'b00;
		`endif
    `endif

    
    reg [7:0] waq;
    
    wire clk_in = (clksel[0] == 1'b0) ? clk0 : clk1;
    wire clk_in_g = (clksel[1] == 1'b0) ? 1'b0 : clk_in;
	
    wire clk_in_d;     

    always @ (posedge clk_in_g)
        waq <= wa;
    
    buf #(1) (clk_in_d, clk_in_g);

    // 2to4 decoder of weq
    wire waq7b_m = ~(waq[7] & we_mode[1]);
    wire waq7_m = ~(waq7b_m & we_mode[1]);
    wire waq7_mg = waq7_m & clk_in_d;
    wire waq7b_mg = waq7b_m & clk_in_d;
    
    wire waq6b_m = ~(waq[6] & we_mode[0]);
    wire waq6_m = ~(waq6b_m & we_mode[0]);
    wire waq6_mg = waq6_m & clk_in_d;
    wire waq6b_mg = waq6b_m & clk_in_d;
    
    assign weq3 = waq7_mg & waq6_mg;
    assign weq2 = waq7_mg & waq6b_mg;
    assign weq1 = waq7b_mg & waq6_mg;
    assign weq0 = waq7b_mg & waq6b_mg;

    // 3to8 decoder of predb
    wire waq4_g = waq[4] & clk_in_d;
    wire waq4b_g = (~waq[4]) & clk_in_d;
    
    wire waq3_g = waq[3] & clk_in_d;
    wire waq3b_g = (~waq[3]) & clk_in_d;
    
    wire waq2_g = waq[2] & clk_in_d;
    wire waq2b_g = (~waq[2]) & clk_in_d;
    
    assign predb[7] = waq4_g & waq3_g & waq2_g;
    assign predb[6] = waq4_g & waq3_g & waq2b_g;
    assign predb[5] = waq4_g & waq3b_g & waq2_g;
    assign predb[4] = waq4_g & waq3b_g & waq2b_g;
    assign predb[3] = waq4b_g & waq3_g & waq2_g;
    assign predb[2] = waq4b_g & waq3_g & waq2b_g;
    assign predb[1] = waq4b_g & waq3b_g & waq2_g;
    assign predb[0] = waq4b_g & waq3b_g & waq2b_g;
    
    //2to4 decoder of preda
    wire waq1_g = waq[1] & clk_in_d;
    wire waq1b_g = (~waq[1]) & clk_in_d;
    
    wire waq0_g = waq[0] & clk_in_d;
    wire waq0b_g = (~waq[0]) & clk_in_d;
    
    assign preda[3] = waq1_g & waq0_g;
    assign preda[2] = waq1_g & waq0b_g;
    assign preda[1] = waq1b_g & waq0_g;
    assign preda[0] = waq1b_g & waq0b_g;
    
    //wa[5]
    assign preda[4] = waq[5];
endmodule

//----------------------------------------------------------------------------
module MUX2S (
    o,
    sel,
    i0,
    i1
);

input        i0;
input        i1;
input        sel;

output        o;

`ifndef CS_SW_SKEL
    assign         o = (sel == 1'b0) ? i0 :
                       (sel == 1'b1) ? i1 : 1'bx;
    specify
        ( i0 =>  o ) = (0,0);                     
        ( i1 =>  o ) = (0,0);                     
        ( sel =>  o ) = (0,0);                                       
    endspecify
`endif

endmodule
//----------------------------------------------------------------------------
//
// module: OSC
//
// description: on-chip oscillator
//
//----------------------------------------------------------------------------


module OSCV1 (
    OSC
);

output OSC;

parameter osc_pd  = 1'b0;
parameter osc_stb = 1'b0;

reg clk;

initial begin
    clk = 1'b0;
    forever #4.76 clk=~clk;
end

assign OSC = osc_pd ? 0 : ( osc_stb ? 0 : clk);

endmodule

module PLLV1 (
    FP_PLL_PDB,  // local signals used to control PLL's power down, low active
    FP_PLL_RST,  // local signals used to control PLL's reset, high active
    fp_cf_clk,
    fp_cf_en,
    fp_cf_in,
    fp_cf_out,
    fp_cf_up,
    fp_cfg_sel,
    PLLCK0       ,  //PLL reference clock0
    PLLCK1       ,  //PLL reference clock1
    FBIN         ,  //feedback clock for deskew mode
    PSEN         ,  // dynamic phase shift enable
    PSCK         ,  // dynamic phase shift clock
    PSDIR        ,  // dynamic phase shift direction
    CO0          ,  //PLL output clock channel 0
    CO1          ,  //PLL output clock channel 1
    CO2          ,  //PLL output clock channel 2
    CO3          ,  //PLL output clock channel 3
    CO4          ,  //PLL output clock channel 4
    CO5          ,  //PLL output clock channel 5
    FBOUT        ,  //PLL feedback clock
    ACTIVECK     ,  //Indicated that which clock is selected now
    CKBAD0       ,  //Indicated PLLCK0 clock is bad
    CKBAD1       ,  //Indicated PLLCK1 clock is bad
    PSDONE       ,  // dynamic phase shift status flag
    PLOCK           //PLL lock status output
`ifdef FM_HACK
    ,CFG_CKSEL
    ,CFG_CK_SWITCH_EN
    ,CFG_SEL_FBPATH
    ,CFG_DIVN
    ,CFG_DIVM
    ,CFG_DIVFB
    ,CFG_LPF
    ,CFG_CPSEL_CR
    ,CFG_CPSEL_FN
    ,CFG_CP_AUTO_ENB
    ,CFG_RST_REG_ENB
    ,CFG_CALIB_EN
    ,CFG_CALIB_RSTN
    ,CFG_CALIB_MANUAL
    ,CFG_CALIB_WIN
    ,CFG_CALIB_DIV
    ,CFG_CALIB_16_32U
    ,CFG_BP_VDOUT
    ,CFG_LKD_MUX
    ,CFG_FORCE_LOCK
    ,CFG_FLDD
    ,CFG_ATEST_EN
    ,CFG_DTEST_EN
    ,CFG_ATEST_SEL
    ,CFG_DTEST_SEL
    ,CFG_VCO_INI_SEL
    ,CFG_LKD_TOL
    ,CFG_LKD_HOLD
    ,CFG_VRSEL
    ,CFG_BK
    ,CFG_SSEN
    ,CFG_SSDIVH
    ,CFG_SSDIVL
    ,CFG_PSSEL
    ,CFG_SSRG
    ,CFG_MKEN0
    ,CFG_MKEN1
    ,CFG_MKEN2
    ,CFG_MKEN3
    ,CFG_MKEN4
    ,CFG_MKEN5
    ,CFG_BPS0
    ,CFG_BPS1
    ,CFG_BPS2
    ,CFG_BPS3
    ,CFG_BPS4
    ,CFG_BPS5
    ,CFG_FRAC
    ,CFG_DIVC0
    ,CFG_DIVC1
    ,CFG_DIVC2
    ,CFG_DIVC3
    ,CFG_DIVC4
    ,CFG_DIVC5
    ,CFG_CO0DLY
    ,CFG_CO1DLY
    ,CFG_CO2DLY
    ,CFG_CO3DLY
    ,CFG_CO4DLY
    ,CFG_CO5DLY
    ,CFG_P0SEL
    ,CFG_P1SEL
    ,CFG_P2SEL
    ,CFG_P3SEL
    ,CFG_P4SEL
    ,CFG_P5SEL
    ,CFG_PFBSEL
    ,CFG_RSTPLL_SEL
    ,CFG_PPDB_SEL
    ,CFG_FP_EN
    ,CFG_LOCK_GATE
`endif
);

//port definition

input         FP_PLL_PDB;
input         FP_PLL_RST;
input         fp_cf_clk;
input         fp_cf_en;
input         fp_cf_in;
output        fp_cf_out;
input         fp_cf_up;
input         fp_cfg_sel;

input         PLLCK0       ;  //PLL reference clock0
input         PLLCK1       ;  //PLL reference clock1
input         FBIN         ;  //feedback clock for deskew mode
input         PSEN         ;  // dynamic phase shift enable
input         PSCK         ;  // dynamic phase shift clock
input         PSDIR        ;  // dynamic phase shift direction


output        CO0          ;  //PLL output clock channel 0
output        CO1          ;  //PLL output clock channel 1
output        CO2          ;  //PLL output clock channel 2
output        CO3          ;  //PLL output clock channel 3
output        CO4          ;  //PLL output clock channel 4
output        CO5          ;  //PLL output clock channel 5
output        FBOUT        ;  //PLL feedback clock output
output        ACTIVECK     ;  //Indicated that which clock is selected now
output        CKBAD0       ;  //Indicated PLLCK0 clock is bad
output        CKBAD1       ;  //Indicated PLLCK1 clock is bad
output        PSDONE       ;  // dynamic phase shift status flag
output        PLOCK        ;  //PLL lock status output

`ifdef FM_HACK
input       CFG_CKSEL        ;
input       CFG_CK_SWITCH_EN ;
input       CFG_SEL_FBPATH   ;
input [7:0] CFG_DIVN         ;
input [7:0] CFG_DIVM         ;
input       CFG_DIVFB        ;
input [2:0] CFG_LPF          ;
input [2:0] CFG_CPSEL_CR     ;
input [6:0] CFG_CPSEL_FN     ;
input       CFG_CP_AUTO_ENB  ;
input       CFG_RST_REG_ENB  ;
input       CFG_CALIB_EN     ;
input       CFG_CALIB_RSTN   ;
input [3:0] CFG_CALIB_MANUAL ;
input [1:0] CFG_CALIB_WIN    ;
input [7:0] CFG_CALIB_DIV    ;
input       CFG_CALIB_16_32U ;
input       CFG_BP_VDOUT     ;
input       CFG_LKD_MUX      ;
input       CFG_FORCE_LOCK   ;
input [1:0] CFG_FLDD         ;
input       CFG_ATEST_EN     ;
input       CFG_DTEST_EN     ;
input       CFG_ATEST_SEL    ;
input       CFG_DTEST_SEL    ;
input       CFG_VCO_INI_SEL  ;
input       CFG_LKD_TOL      ;
input       CFG_LKD_HOLD     ;
input [1:0] CFG_VRSEL        ;
input [3:0] CFG_BK           ;
input       CFG_SSEN         ;
input [1:0] CFG_SSDIVH       ;
input [7:0] CFG_SSDIVL       ;
input [5:0] CFG_PSSEL        ;
input [1:0] CFG_SSRG         ;
input       CFG_MKEN0        ;
input       CFG_MKEN1        ;
input       CFG_MKEN2        ;
input       CFG_MKEN3        ;
input       CFG_MKEN4        ;
input       CFG_MKEN5        ;
input       CFG_BPS0         ;
input       CFG_BPS1         ;
input       CFG_BPS2         ;
input       CFG_BPS3         ;
input       CFG_BPS4         ;
input       CFG_BPS5         ;
input [2:0] CFG_FRAC         ;
input [7:0] CFG_DIVC0        ;
input [7:0] CFG_DIVC1        ;
input [7:0] CFG_DIVC2        ;
input [7:0] CFG_DIVC3        ;
input [7:0] CFG_DIVC4        ;
input [7:0] CFG_DIVC5        ;
input [7:0] CFG_CO0DLY       ;
input [7:0] CFG_CO1DLY       ;
input [7:0] CFG_CO2DLY       ;
input [7:0] CFG_CO3DLY       ;
input [7:0] CFG_CO4DLY       ;
input [7:0] CFG_CO5DLY       ;
input [2:0] CFG_P0SEL        ;
input [2:0] CFG_P1SEL        ;
input [2:0] CFG_P2SEL        ;
input [2:0] CFG_P3SEL        ;
input [2:0] CFG_P4SEL        ;
input [2:0] CFG_P5SEL        ;
input [2:0] CFG_PFBSEL       ;
input [1:0] CFG_RSTPLL_SEL   ;
input [1:0] CFG_PPDB_SEL     ;
input       CFG_FP_EN        ;
input       CFG_LOCK_GATE    ;
`else
parameter    pll_sel = "auto"; //default: "auto", can be "0", "1", "2" or "3".

parameter    CFG_CKSEL        = 1'b0;  //PLL reference clk sel when ck_switch off
parameter    CFG_CK_SWITCH_EN = 1'b0;  // Input clock automatic selection enable 0:manual select  (default) 1:automatic select
parameter    CFG_SEL_FBPATH   = 1'b0;  //select the feedback signal to PFD
parameter    CFG_DIVN         = 8'b0;  //input divider control
parameter    CFG_DIVM         = 8'b0;  //loop divider control
parameter    CFG_DIVFB        = 1'b0;  //internal feedback clock of VCO control 1:bypass. 0:divide by 2
parameter    CFG_LPF          = 3'b0;  //loop filter resistance value adjustment
parameter    CFG_CPSEL_CR     = 3'b0;  //select CP current,coarse tune
parameter    CFG_CPSEL_FN     = 7'b0;  //select CP current,fine tune
parameter    CFG_CP_AUTO_ENB  = 1'b0;  //cp current control sel
parameter    CFG_RST_REG_ENB  = 1'b0;  //internal regulator por signal control
parameter    CFG_CALIB_EN     = 1'b0;  // vco calibration enable 
parameter    CFG_CALIB_RSTN   = 1'b0;  // vco calibration reset
parameter    CFG_CALIB_MANUAL = 4'b0;  // vco calibration manual mode
parameter    CFG_CALIB_WIN    = 2'b0;  // vco calibration vc monitor voltage window sel
parameter    CFG_CALIB_DIV    = 8'b0;  // vco calibration clock divider setting
parameter    CFG_CALIB_16_32U = 1'b0;  // vco calibration time sel
parameter    CFG_BP_VDOUT     = 1'b0;  //bypass dvdd(core) to vddd
parameter    CFG_LKD_MUX      = 1'b0;  //lock detector ref clk sel 0: feedback clk 1:reference clk
parameter    CFG_FORCE_LOCK   = 1'b0;  //force PLOCK signal to high
parameter    CFG_FLDD         = 2'b0;  //lock detector range select
parameter    CFG_ATEST_EN     = 1'b0;  //test control enable for analog test 
parameter    CFG_DTEST_EN     = 1'b0;  //test control enable for digital test 
parameter    CFG_ATEST_SEL    = 1'b0;  //analog test select
parameter    CFG_DTEST_SEL    = 1'b0;  //digital test select
parameter    CFG_VCO_INI_SEL  = 1'b0;  //vco initial phase align control
parameter    CFG_LKD_TOL      = 1'b0;  //Lock Detector tolerance (TBD)
parameter    CFG_LKD_HOLD     = 1'b0;  // Lock Detector hold number (TBD) 
parameter    CFG_VRSEL        = 2'b0;  //select the reference voltage for regulator
parameter    CFG_BK           = 4'b0;  //Back up register 
parameter    CFG_SSEN         = 1'b0;  //Spread spectrum function enable 0:don't use SSCG function  (default) 1:enable
parameter    CFG_SSDIVH       = 2'b0;  //Spread frequency-divider 1 control, range within[1,16] divider value NH=SSDIVH<3:0>+1
parameter    CFG_SSDIVL       = 8'b0;  //Spread frequency-divider 2 control, range within[1,256] divider value NH=SSDIVL<7:0>+1
parameter    CFG_PSSEL        = 6'b0;  // dynamic phase shift channel sel
parameter    CFG_SSRG         = 2'b0;  //Spread ratio select (TBD)
parameter    CFG_MKEN0        = 1'b0;  //output enable for channel 0
parameter    CFG_MKEN1        = 1'b0;  //output enable for channel 1
parameter    CFG_MKEN2        = 1'b0;  //output enable for channel 2
parameter    CFG_MKEN3        = 1'b0;  //output enable for channel 3
parameter    CFG_MKEN4        = 1'b0;  //output enable for channel 4
parameter    CFG_MKEN5        = 1'b0;  //output enable for channel 5
parameter    CFG_BPS0         = 1'b0;  //bypass output of channel 0
parameter    CFG_BPS1         = 1'b0;  //bypass output of channel 1
parameter    CFG_BPS2         = 1'b0;  //bypass output of channel 2
parameter    CFG_BPS3         = 1'b0;  //bypass output of channel 3
parameter    CFG_BPS4         = 1'b0;  //bypass output of channel 4
parameter    CFG_BPS5         = 1'b0;  //bypass output of channel 5
parameter    CFG_FRAC         = 3'b0;  //Frac-divider setting
parameter    CFG_DIVC0        = 8'b0;  //output divider control for channel 0
parameter    CFG_DIVC1        = 8'b0;  //output divider control for channel 1
parameter    CFG_DIVC2        = 8'b0;  //output divider control for channel 2
parameter    CFG_DIVC3        = 8'b0;  //output divider control for channel 3
parameter    CFG_DIVC4        = 8'b0;  //output divider control for channel 4
parameter    CFG_DIVC5        = 8'b0;  //output divider control for channel 5
parameter    CFG_CO0DLY       = 8'b0;  //channel 0 coarse delay control
parameter    CFG_CO1DLY       = 8'b0;  //channel 1 coarse delay control
parameter    CFG_CO2DLY       = 8'b0;  //channel 2 coarse delay control
parameter    CFG_CO3DLY       = 8'b0;  //channel 3 coarse delay control
parameter    CFG_CO4DLY       = 8'b0;  //channel 4 coarse delay control
parameter    CFG_CO5DLY       = 8'b0;  //channel 5 coarse delay control
parameter    CFG_P0SEL        = 3'b0;  //select phase for channel 0
parameter    CFG_P1SEL        = 3'b0;  //select phase for channel 1
parameter    CFG_P2SEL        = 3'b0;  //select phase for channel 2
parameter    CFG_P3SEL        = 3'b0;  //select phase for channel 3
parameter    CFG_P4SEL        = 3'b0;  //select phase for channel 4
parameter    CFG_P5SEL        = 3'b0;  //select phase for channel 5
parameter    CFG_PFBSEL       = 3'b0;  //select phase for feedback clock

parameter    CFG_RSTPLL_SEL   = 2'b0;
parameter    CFG_PPDB_SEL     = 2'b0; //Controlled by Fabric.
parameter    CFG_FP_EN        = 1'b0;

parameter    CFG_LOCK_GATE    = 1'b0;
`endif

wire         PDB          ;  //power-down mode control
wire         RSTPLL       ;  //reset PLL control

wire  [2:0]  FP_LPF      ;
wire  [2:0]  FP_CPSEL_CR ;
wire  [7:0]  FP_DIVN     ;
wire  [7:0]  FP_DIVM     ;
wire  [7:0]  FP_DIVC5    ;
wire  [7:0]  FP_DIVC4    ;
wire  [7:0]  FP_DIVC3    ;
wire  [7:0]  FP_DIVC2    ;
wire  [7:0]  FP_DIVC1    ;
wire         FP_MKEN5    ;
wire         FP_MKEN4    ;
wire         FP_MKEN3    ;
wire         FP_MKEN2    ;
wire         FP_MKEN1    ;
wire         FP_MKEN0    ;
wire  [2:0]  FP_FRAC     ;
wire  [7:0]  FP_DIVC0    ;
wire         FP_DIVFB    ;

reg por;
initial begin
    por = 1'b0;
    #5;
    por = 1'b1;
end

reg [79:0] cfg_dyn_dff;
reg [79:0] cfg_dyn_lat;

always@(posedge fp_cf_clk or negedge por)
begin
    if(~por)
        cfg_dyn_dff <= 0;
    else if(fp_cf_en)
        cfg_dyn_dff <= {cfg_dyn_dff,fp_cf_in};
end

assign fp_cf_out = fp_cf_en & cfg_dyn_dff[79];

always@(posedge fp_cf_up or negedge por)
begin
    if(~por)
        cfg_dyn_lat <= 0;
    else
        cfg_dyn_lat <= cfg_dyn_dff;
end

assign {FP_LPF[2:0], 
        FP_CPSEL_CR[2:0], 
        FP_DIVN[7:0], 
        FP_DIVM[7:0], 
        FP_DIVC5[7:0], 
        FP_DIVC4[7:0], 
        FP_DIVC3[7:0], 
        FP_DIVC2[7:0], 
        FP_DIVC1[7:0], 
        FP_MKEN5, 
        FP_MKEN4, 
        FP_MKEN3, 
        FP_MKEN2, 
        FP_MKEN1, 
        FP_MKEN0, 
        FP_FRAC[2:0], 
        FP_DIVC0[7:0], 
        FP_DIVFB
       } = cfg_dyn_lat;

assign RSTPLL = CFG_RSTPLL_SEL[1:0] == 2'b11 ? FP_PLL_RST   : //Controlled by Fabric.
                CFG_RSTPLL_SEL[1:0] == 2'b10 ? 1'b1         : //control by reg
                CFG_RSTPLL_SEL[1:0] == 2'b01 ? 1'b0         : //non-reset
                                               1'b1         ; //reset

assign PDB   = CFG_PPDB_SEL[1:0] == 2'b11 ? FP_PLL_PDB   : //Controlled by Fabric.
               CFG_PPDB_SEL[1:0] == 2'b10 ? 1'b1         : //control by reg
               CFG_PPDB_SEL[1:0] == 2'b01 ? 1'b1         : //always on
                                            1'b0         ; //always off

wire         CKSEL        = CFG_CKSEL        ;
wire         CK_SWITCH_EN = CFG_CK_SWITCH_EN ;
wire         SEL_FBPATH   = CFG_SEL_FBPATH   ;
wire  [6:0]  CPSEL_FN     = CFG_CPSEL_FN     ;
wire         CP_AUTO_ENB  = CFG_CP_AUTO_ENB  ;
wire         RST_REG_ENB  = CFG_RST_REG_ENB  ;
wire         CALIB_EN     = CFG_CALIB_EN     ;
wire         CALIB_RSTN   = CFG_CALIB_RSTN   ;
wire  [3:0]  CALIB_MANUAL = CFG_CALIB_MANUAL ;
wire  [1:0]  CALIB_WIN    = CFG_CALIB_WIN    ;
wire  [7:0]  CALIB_DIV    = CFG_CALIB_DIV    ;
wire         CALIB_16_32U = CFG_CALIB_16_32U ;
wire         BP_VDOUT     = CFG_BP_VDOUT     ;
wire         LKD_MUX      = CFG_LKD_MUX      ;
wire         FORCE_LOCK   = CFG_FORCE_LOCK   ;
wire  [1:0]  FLDD         = CFG_FLDD         ;
wire         ATEST_EN     = CFG_ATEST_EN     ;
wire         DTEST_EN     = CFG_DTEST_EN     ;
wire         ATEST_SEL    = CFG_ATEST_SEL    ;
wire         DTEST_SEL    = CFG_DTEST_SEL    ;
wire         VCO_INI_SEL  = CFG_VCO_INI_SEL  ;
wire         LKD_TOL      = CFG_LKD_TOL      ;
wire         LKD_HOLD     = CFG_LKD_HOLD     ;
wire  [1:0]  VRSEL        = CFG_VRSEL        ;
wire  [3:0]  BK           = CFG_BK           ;
wire         SSEN         = CFG_SSEN         ;
wire  [1:0]  SSDIVH       = CFG_SSDIVH       ;
wire  [7:0]  SSDIVL       = CFG_SSDIVL       ;
wire  [5:0]  PSSEL        = CFG_PSSEL        ;
wire  [1:0]  SSRG         = CFG_SSRG         ;
wire         BPS0         = CFG_BPS0         ;
wire         BPS1         = CFG_BPS1         ;
wire         BPS2         = CFG_BPS2         ;
wire         BPS3         = CFG_BPS3         ;
wire         BPS4         = CFG_BPS4         ;
wire         BPS5         = CFG_BPS5         ;
wire  [7:0]  CO0DLY       = CFG_CO0DLY       ;
wire  [7:0]  CO1DLY       = CFG_CO1DLY       ;
wire  [7:0]  CO2DLY       = CFG_CO2DLY       ;
wire  [7:0]  CO3DLY       = CFG_CO3DLY       ;
wire  [7:0]  CO4DLY       = CFG_CO4DLY       ;
wire  [7:0]  CO5DLY       = CFG_CO5DLY       ;
wire  [2:0]  P0SEL        = CFG_P0SEL        ;
wire  [2:0]  P1SEL        = CFG_P1SEL        ;
wire  [2:0]  P2SEL        = CFG_P2SEL        ;
wire  [2:0]  P3SEL        = CFG_P3SEL        ;
wire  [2:0]  P4SEL        = CFG_P4SEL        ;
wire  [2:0]  P5SEL        = CFG_P5SEL        ;
wire  [2:0]  PFBSEL       = CFG_PFBSEL       ;

wire  [2:0]  LPF          = CFG_FP_EN & fp_cfg_sel ? FP_LPF[2:0]      : CFG_LPF[2:0]      ;
wire  [2:0]  CPSEL_CR     = CFG_FP_EN & fp_cfg_sel ? FP_CPSEL_CR[2:0] : CFG_CPSEL_CR[2:0] ;
wire  [7:0]  DIVN         = CFG_FP_EN & fp_cfg_sel ? FP_DIVN[7:0]     : CFG_DIVN[7:0]     ;
wire  [7:0]  DIVM         = CFG_FP_EN & fp_cfg_sel ? FP_DIVM[7:0]     : CFG_DIVM[7:0]     ;
wire  [7:0]  DIVC5        = CFG_FP_EN & fp_cfg_sel ? FP_DIVC5[7:0]    : CFG_DIVC5[7:0]    ;
wire  [7:0]  DIVC4        = CFG_FP_EN & fp_cfg_sel ? FP_DIVC4[7:0]    : CFG_DIVC4[7:0]    ;
wire  [7:0]  DIVC3        = CFG_FP_EN & fp_cfg_sel ? FP_DIVC3[7:0]    : CFG_DIVC3[7:0]    ;
wire  [7:0]  DIVC2        = CFG_FP_EN & fp_cfg_sel ? FP_DIVC2[7:0]    : CFG_DIVC2[7:0]    ;
wire  [7:0]  DIVC1        = CFG_FP_EN & fp_cfg_sel ? FP_DIVC1[7:0]    : CFG_DIVC1[7:0]    ;
wire         MKEN5        = CFG_FP_EN & fp_cfg_sel ? FP_MKEN5         : CFG_MKEN5         ;
wire         MKEN4        = CFG_FP_EN & fp_cfg_sel ? FP_MKEN4         : CFG_MKEN4         ;
wire         MKEN3        = CFG_FP_EN & fp_cfg_sel ? FP_MKEN3         : CFG_MKEN3         ;
wire         MKEN2        = CFG_FP_EN & fp_cfg_sel ? FP_MKEN2         : CFG_MKEN2         ;
wire         MKEN1        = CFG_FP_EN & fp_cfg_sel ? FP_MKEN1         : CFG_MKEN1         ;
wire         MKEN0        = CFG_FP_EN & fp_cfg_sel ? FP_MKEN0         : CFG_MKEN0         ;
wire  [2:0]  FRAC         = CFG_FP_EN & fp_cfg_sel ? FP_FRAC[2:0]     : CFG_FRAC[2:0]     ;
wire  [7:0]  DIVC0        = CFG_FP_EN & fp_cfg_sel ? FP_DIVC0[7:0]    : CFG_DIVC0[7:0]    ;
wire         DIVFB        = CFG_FP_EN & fp_cfg_sel ? FP_DIVFB         : CFG_DIVFB         ;

supply1         VDDIO        ;  //io power supply for regulator  
supply0         VSSIO        ;  //io ground for regulator
supply1         DVDD         ;  //digital power supply
supply0         DVSS         ;  //digital ground
supply0         AVSS_VCO     ;  //VCO ground
supply0         AVSS         ;  //analog ground
supply1         VREF         ;  //reference voltage for regulator

wire [1:0] dangling;

PLL_TOP PLL_TOP (
	.VDDIO		(VDDIO),
	.VSSIO		(VSSIO),
	.DVDD		(DVDD),
	.DVSS		(DVSS),
	.AVSS_VCO	(AVSS_VCO),
	.AVSS		(AVSS),
	.PLLCK0		(PLLCK0),
	.PLLCK1		(PLLCK1),
	.FBIN		(FBIN),
	.VREF		(VREF),
	.CKSEL		(CKSEL),
	.CK_SWITCH_EN	(CK_SWITCH_EN),
	.PDB		(PDB),
	.RSTPLL		(RSTPLL),
	.SEL_FBPATH	(SEL_FBPATH),
	.DIVN		(DIVN[7:0]),
	.DIVM		(DIVM[7:0]),
	.DIVFB		(DIVFB),
	.LPF		(LPF[2:0]),
	.CPSEL_CR	(CPSEL_CR[2:0]),
	.CPSEL_FN	(CPSEL_FN[6:0]),
	.CP_AUTO_ENB	(CP_AUTO_ENB),
	.RST_REG_ENB	(RST_REG_ENB),
	.CALIB_EN	(CALIB_EN),
	.CALIB_RSTN	(CALIB_RSTN),
	.CALIB_MANUAL	(CALIB_MANUAL[3:0]),
	.CALIB_WIN	(CALIB_WIN[1:0]),
	.CALIB_DIV	(CALIB_DIV[7:0]),
	.CALIB_16_32U	(CALIB_16_32U),
	.BP_VDOUT	(BP_VDOUT),
	.LKD_MUX	(LKD_MUX),
	.FORCE_LOCK	(FORCE_LOCK),
	.FLDD		(FLDD[1:0]),
	.ATEST_EN	(ATEST_EN),
	.DTEST_EN	(DTEST_EN),
	.ATEST_SEL	(ATEST_SEL),
	.DTEST_SEL	(DTEST_SEL),
	.VCO_INI_SEL	(VCO_INI_SEL),
	.LKD_TOL	(LKD_TOL),
	.LKD_HOLD	(LKD_HOLD),
	.VRSEL		(VRSEL[1:0]),
	.BK		(BK[3:0]),
	.SSEN		(SSEN),
	.SSDIVH		(SSDIVH[1:0]),
	.SSDIVL		(SSDIVL[7:0]),
	.SSRG		(SSRG[1:0]),
	.PSEN		(PSEN),
	.PSCK		(PSCK),
	.PSDIR		(PSDIR),
	.PSSEL		(PSSEL[5:0]),
	.MKEN0		(MKEN0),
	.MKEN1		(MKEN1),
	.MKEN2		(MKEN2),
	.MKEN3		(MKEN3),
	.MKEN4		(MKEN4),
	.MKEN5		(MKEN5),
	.BPS0		(BPS0),
	.BPS1		(BPS1),
	.BPS2		(BPS2),
	.BPS3		(BPS3),
	.BPS4		(BPS4),
	.BPS5		(BPS5),
	.FRAC		(FRAC[2:0]),
	.DIVC0		(DIVC0[7:0]),
	.DIVC1		(DIVC1[7:0]),
	.DIVC2		(DIVC2[7:0]),
	.DIVC3		(DIVC3[7:0]),
	.DIVC4		(DIVC4[7:0]),
	.DIVC5		(DIVC5[7:0]),
	.CO0DLY		(CO0DLY[7:0]),
	.CO1DLY		(CO1DLY[7:0]),
	.CO2DLY		(CO2DLY[7:0]),
	.CO3DLY		(CO3DLY[7:0]),
	.CO4DLY		(CO4DLY[7:0]),
	.CO5DLY		(CO5DLY[7:0]),
	.P0SEL		(P0SEL[2:0]),
	.P1SEL		(P1SEL[2:0]),
	.P2SEL		(P2SEL[2:0]),
	.P3SEL		(P3SEL[2:0]),
	.P4SEL		(P4SEL[2:0]),
	.P5SEL		(P5SEL[2:0]),
	.PFBSEL		(PFBSEL[2:0]),

	.CO0		(CO0_t),
	.CO1		(CO1_t),
	.CO2		(CO2_t),
	.CO3		(CO3_t),
	.CO4		(CO4_t),
	.CO5		(CO5_t),
	.FBOUT		(FBOUT_t),
	.ACTIVECK	(ACTIVECK),
	.CKBAD0		(CKBAD0),
	.CKBAD1		(CKBAD1),
	.PSDONE		(PSDONE),
	.PLOCK		(PLOCK),
	.ATEST_PLL	(dangling[0]),
	.DTEST_PLL	(dangling[1]) 
);

co_lock_gate u0_gate (.TE(CFG_LOCK_GATE), .E(PLOCK), .CP(CO0_t), .Q(CO0));
co_lock_gate u1_gate (.TE(CFG_LOCK_GATE), .E(PLOCK), .CP(CO1_t), .Q(CO1));
co_lock_gate u2_gate (.TE(CFG_LOCK_GATE), .E(PLOCK), .CP(CO2_t), .Q(CO2));
co_lock_gate u3_gate (.TE(CFG_LOCK_GATE), .E(PLOCK), .CP(CO3_t), .Q(CO3));
co_lock_gate u4_gate (.TE(CFG_LOCK_GATE), .E(PLOCK), .CP(CO4_t), .Q(CO4));
co_lock_gate u5_gate (.TE(CFG_LOCK_GATE), .E(PLOCK), .CP(CO5_t), .Q(CO5));
co_lock_gate fb_gate (.TE(vcc),           .E(vcc),   .CP(FBOUT_t), .Q(FBOUT));
supply1_guts V (.vcc(vcc));
 
endmodule

//----------------------------------------------------------------------------
//
// module: REG2CKSR
//
// description: 1 bit register or latch with "sr" to preset value
//		to use as latch, hold mclk_b=0 (master stage transparent)
//		Two clock inputs, config-mux selectable
// config:      PRESET, CLKSRSEL
//
//----------------------------------------------------------------------------
module REG2CKSR (
    qx,
    di,
    sr0,
    sr1,
    mclk0b,
    sclk0,
    mclk1b,
    sclk1
`ifdef FM_HACK
	,PRESET
	,CLKSRSEL
`endif
);

output        qx;

input         di;
input         sr0, sr1;
input         mclk0b;
input         sclk0;
input         mclk1b;
input         sclk1;


`ifdef CS_FORMALPRO_HACK
   wire        PRESET;
   wire        CLKSRSEL;
`else
     `ifdef  SIMULATION
          reg       PRESET   = 1'b0;
          reg       CLKSRSEL = 1'b0;
     `else
		`ifdef FM_HACK
	        input PRESET;
	        input CLKSRSEL;
		`else
	        parameter PRESET   = 1'b0;
	        parameter CLKSRSEL = 1'b0;
		`endif
     `endif
`endif

wire            mclkb;
wire            sclk;
   reg          qx_reg;
   reg          mout;

`ifndef CS_SW_SKEL



   assign    mclkb = (CLKSRSEL == 1'b1) ? mclk1b : mclk0b;
   assign    sclk   = (CLKSRSEL == 1'b1) ? sclk1   : sclk0;
 
   wire    a_sr = (CLKSRSEL == 1'b1) ? sr1: sr0;
   wire    rst_ =  a_sr || (PRESET == 1'b1);
   wire    set  = ~a_sr && (PRESET == 1'b1);    
  
   always @(*) begin
       if (rst_ == 1'b0) begin
           mout <= 1;
       end else if (set) begin
           mout <= 0;
       end else if (mclkb == 0) begin
           mout <= ~di;
       end else if (mclkb == 1) begin
           mout <= mout;
       end else
           mout <= 1'bx;
   end

   initial qx_reg = 1'b0;
   
   always @(*) begin
       if (rst_ == 1'b0) begin
           qx_reg <= 1;
       end else if (set) begin
           qx_reg <= 0;
       end else if (sclk == 1) begin
           qx_reg <= mout;
       end else if (sclk == 0) begin
           qx_reg <= qx_reg;
       end else
           qx_reg <= 1'bx;
   end 
   
   assign qx = ~qx_reg;

    specify
        (posedge sclk0 => ( qx  +: di) ) = (0, 0) ;
        (posedge sclk1 => ( qx  +: di) ) = (0, 0) ;
              
        $setuphold(posedge sclk, di, 0, 0);
        $recrem(a_sr, posedge sclk,  0, 0);
        
     endspecify
   

`endif

endmodule

module SOC_SLAVE_BUS(
    fpinf_write,
    fpinf_addr,
    fpinf_req,
    fpinf_gnt,
    fpinf_wdata,
    fpinf_rdata,
    fp_rcfg_req,
    rst_fpinf_n
);

output             fpinf_write;
output   [7:0]     fpinf_addr;
output             fpinf_req;
input              fpinf_gnt;
output   [15:0]    fpinf_wdata;
input    [15:0]    fpinf_rdata;
input              fp_rcfg_req;
input              rst_fpinf_n;

parameter fp_rcfg_en     = 1'b0;
parameter fp_recfg_addr  = 24'h0;

endmodule

//----------------------------------------------------------------------------
//
// module: SUPPLY 0
//
// description: GND Cell
//
//----------------------------------------------------------------------------
module supply0_guts (
            gnd
	     );

    output		gnd;

assign gnd = 0;
endmodule
//----------------------------------------------------------------------------
//
// module: SUPPLY 1
//
// description: vcc Cell
//
//----------------------------------------------------------------------------
module supply1_guts (
            vcc
         );

    output      vcc;

assign vcc = 1;
endmodule

module UPDATE(
	update,
	update_,
	align_user,
	geclk0
	`ifdef FM_HACK
	,CFG_UP_SEL
	`endif
	);
output	update,update_;
input	align_user;
input	geclk0;
`ifdef FM_HACK
input	[6:0]	CFG_UP_SEL;
`else
parameter	[6:0]	CFG_UP_SEL=7'b000_0000;
`endif
`ifndef FM_HACK
reg usermode;
wire GSR;
glbsr inst( .GSR( GSR )) ;

initial begin
    usermode = 1'b0;
	@(posedge GSR);
	usermode = 1'b1;
end
`else
wire usermode = 1'b1;
`endif
wire usermode_b = ~usermode;
//align user logic
iob_dff a0(.q(align_a),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(1'b1),.d(align_user));
iob_dff a1(.q(align_b),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(1'b1),.d(align_a));
iob_dff a2(.q(align_cn),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(1'b1),.d(align_b));
wire align_n = !(align_b & ~align_cn);
/////////////////////////////
//update shift register loop
IO_MUX2S1 m7(.o(d0),.in0(q3),.in1(q7),.SEL(CFG_UP_SEL[6]));
IO_MUX2S1 m6(.o(d7),.in0(q6),.in1(q4),.SEL(CFG_UP_SEL[3]));
IO_MUX2S1 m5(.o(d6),.in0(q5),.in1(q4),.SEL(CFG_UP_SEL[4]));
IO_MUX2S1 m4(.o(d5),.in0(1'b1),.in1(q4),.SEL(CFG_UP_SEL[5]));
IO_MUX2S1 m3(.o(d4),.in0(1'b1),.in1(q3),.SEL(CFG_UP_SEL[6]));
IO_MUX2S1 m2(.o(d3),.in0(q2),.in1(q0),.SEL(CFG_UP_SEL[0]));
IO_MUX2S1 m1(.o(d2),.in0(q1),.in1(q0),.SEL(CFG_UP_SEL[1]));
IO_MUX2S1 m0(.o(d1),.in0(1'b1),.in1(q0),.SEL(CFG_UP_SEL[2]));
iob_dff u0(.q(q0),.clk(geclk0),.rst(1'b0),.set_(usermode),.en(align_n),.d(d0));
iob_dff u1(.q(q1),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d1));
iob_dff u2(.q(q2),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d2));
iob_dff u3(.q(q3),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d3));
iob_dff u4(.q(q4),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d4));
iob_dff u5(.q(q5),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d5));
iob_dff u6(.q(q6),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d6));
iob_dff u7(.q(q7),.clk(geclk0),.rst(usermode_b),.set_(1'b1),.en(align_n),.d(d7));
////////////////////////////
assign update  = d0;
assign update_ = ~d0;
endmodule
module cts_dffrs(D,CK,Q,QB,SETN,RSTN);
input D,CK;
output Q,QB;
input SETN,RSTN;
reg Q;

assign QB=~Q;

always @(posedge CK or negedge SETN or negedge RSTN) begin
    if(RSTN==0)
        Q<=0;
    else if(SETN==0)
        Q<=1;
    else
        Q<=D;
end
endmodule



module SDLLV1(
     DQS
    ,DQS_O
    ,SOF
    ,SUF
    ,CLKUP
    ,DCTLIN
    ,START_S
    ,DOFF
    ,FBSEL
    ,SSEL
    ,BK
);

//input
input            DQS         ;
input            CLKUP       ;
input    [9:0]   DCTLIN      ;

//output
output            DQS_O      ;
output            SOF        ;
output            SUF        ;

input            START_S     ;
input    [4:0]   DOFF        ;
input    [1:0]   FBSEL       ;
input    [3:0]   SSEL        ;
input    [1:0]   BK          ;

supply0 VSS;
supply1 VDD;

SDLL_TOP sdll(
     .DVDD          ( VDD     )
    ,.DVSS          ( VSS     )
    ,.DVDDL         ( VDD     )
    ,.DVSSL         ( VSS     )
    ,.DQS           ( DQS     )
    ,.DQS_O         ( DQS_O   )
    ,.SOF           ( SOF     )
    ,.SUF           ( SUF     )
    ,.DCTLIN        ( DCTLIN  )
    ,.CLKUP         ( CLKUP   )
    ,.DOFF          ( DOFF    )
    ,.START_S       ( START_S )
    ,.FBSEL         ( FBSEL   )
    ,.SSEL          ( SSEL    )
    ,.BK            ( BK      )
);

endmodule

module MDLLV1(
     DLLCK
    ,CKOUT
    ,DCTLO
    ,CLKUP
    ,DLOCK
    ,FAIL
    ,OF
    ,UF
    ,DTEST
    ,START
    ,FBSEL
    ,MSEL
    ,DR
    ,DTEST_EN
    ,DTEST_SEL
    ,BK
);
    
//input
input            DLLCK      ;

//output
output          CKOUT       ;
output  [9:0]   DCTLO       ;
output          CLKUP       ;
output          DLOCK       ;
output          FAIL        ;
output          OF          ;
output          UF          ;
output          DTEST       ;

input           START       ;
input   [1:0]   FBSEL       ;
input   [3:0]   MSEL        ;
input           DR          ;
input           DTEST_EN    ;
input   [1:0]   DTEST_SEL   ;
input   [3:0]   BK          ;

supply0 VSS;
supply1 VDD;

MDLL_TOP mdll(
     .DVDD          ( VDD       )
    ,.DVSS          ( VSS       )
    ,.DVDDL         ( VDD       )
    ,.DVSSL         ( VSS       )
    ,.DLLCK         ( DLLCK     )
    ,.CKOUT         ( CKOUT     )
    ,.DCTLO         ( DCTLO     )
    ,.CLKUP         ( CLKUP     )
    ,.DLOCK         ( DLOCK     )
    ,.FAIL          ( FAIL      )
    ,.OF            ( OF        )
    ,.UF            ( UF        )
    ,.DTEST         ( DTEST     )
    ,.START         ( START     )
    ,.FBSEL         ( FBSEL     )
    ,.MSEL          ( MSEL      )
    ,.DR            ( DR        )
    ,.DTEST_EN      ( DTEST_EN  )
    ,.DTEST_SEL     ( DTEST_SEL )
    ,.BK            ( BK        )
);

endmodule



///////////////////////////////////////////////////////////////
// Verilog behavioral model of MDLL (master delay line loop) //
//                                                           //
// Version: 1.0                                              //
// Date:  Jul 18, 2014                                       //
// purpose: for logic behavioral simulation.                 //
// Creator: CME      					     //
// Author:  Zgsu                                             //
// Update information:                                       //
// version 1.0 : basic version                               //   
//                                                           //
///////////////////////////////////////////////////////////////

`timescale 1ns/1ps
module MDLL_TOP(
                   DVDD		,
                   DVSS		,
                   DVDDL	,
                   DVSSL	,
                   DLLCK	,
                   CKOUT	,
                   DCTLO	,
                   CLKUP	,
                   DLOCK	,
                   FAIL		,
                   OF		,
                   UF		,
                   DTEST	,
                   START	,
                   FBSEL	,
                   MSEL		,
                   DR		,
                   DTEST_EN	,
                   DTEST_SEL	,
                   BK
  );

//parameters definition

parameter MAX_INPUT_PERIOD  = 20;	// input range    : 50MHZ-667MHz    
parameter MIN_INPUT_PERIOD  = 1.5;	//   
parameter LOCK_TIME         = 200;	// max lock time=100*INPUT_PERIOD 
    
//port definition

//input
input		DVDD		;  // digital power, share to core power
input		DVSS		;  // digital ground, share to core ground
input		DVDDL		;  // DCDL power, share to core power
input		DVSSL		;  // DCDL ground, share to core ground
input		DLLCK		;  // MDLL reference clock
input		START		;  // MDLL start to work(default:0)
input	[1:0]	FBSEL		;  // how many stages of delay chain to be used.(default:00)
input	[3:0]	MSEL		;  // CKOUT phase select, the phase depend on the FBSEL.(default:0000)
input		DR		;  // divide ratio between the internal controller clock and the input clock.(deault:0)
input		DTEST_EN	;  // DTEST enable.(default:0)
input	[1:0]	DTEST_SEL	;  // DTEST source select
input	[3:0]	BK		;  // BK[3] is minimum delay enable,BK[2:0] for backup.(default:0000)

//output
output		CKOUT		;  // MDLL output clock
output	[9:0]	DCTLO		;  // digital control bits to SDLL
output		CLKUP		;  // synchronous clock with DCTLO, rising edge triggered
output		DLOCK		;  // MDLL lock status indication. 0:no lock, 1:locked
output		FAIL		;  // MDLL failed to lock. 0:normal work, 1:failed
output		OF		;  // MDLL control bits overflow. 0:normal work, 1:overflow
output		UF		;  // MDLL control bits underflow. 0:normal work, 1:underflow
output		DTEST		;  // digital signal test


endmodule
//////////////////////////////////////////////////////////////
// Verilog behavioral model of SDLL (slave delay line loop) //
//                                                          //
// Version: 1.1                                             //
// Date:  Sep 04, 2014                                      //
// purpose: for logic behavioral simulation.                //
// Creator: CME                                             //
// Author:  Zgsu                                            //
// Update information:                                      //
// version 1.0 : basic version                              //   
//         1.1 : update DOFF[3:0] to DOFF[4:0]              //   
//             : add SOF and SUF output pin                 //   
//                                                          //
//////////////////////////////////////////////////////////////

`timescale 1ns/1ps
module SDLL_TOP(
                   DVDD		,
                   DVSS		,
                   DVDDL	,
                   DVSSL	,
                   DQS		,
                   DQS_O	,
                   SOF		,
                   SUF		,
                   DCTLIN	,
                   CLKUP	,
                   DOFF		,
                   START_S	,
                   FBSEL	,
                   SSEL		,
                   BK
  );

//parameters definition

parameter MAX_INPUT_PERIOD  = 20;	// input range    : 50MHZ-667MHz    
parameter MIN_INPUT_PERIOD  = 1.5;	//   
    
//port definition

//input
input		DVDD		;  // digital power, share to core power
input		DVSS		;  // digital ground, share to core ground
input		DVDDL		;  // DCDL power, share to core power
input		DVSSL		;  // DCDL ground, share to core ground
input		DQS		;  // DQS clock, input to SDLL
input		START_S		;  // SDLL start to work(default:0)
input	[9:0]	DCTLIN		;  // digital control bits from MDLL
input		CLKUP		;  // synchronous clock with DCTLIN, rising edge triggered
input	[4:0]	DOFF		;  // delay offset control.(default:00000)
input	[1:0]	FBSEL		;  // how many stages of delay chain to be used.(default:00)
input	[3:0]	SSEL		;  // DQS_O phase select, the phase depend on the FBSEL.(default:0000)
input	[1:0]	BK		;  // BK[1] is minimum delay enable,BK[0] for backup.(default:00)

//output
output		DQS_O		;  // SDLL output clock
output		SOF		;  // SDLL overflow indication
output		SUF		;  // SDLL underflow indication


endmodule
module DNT_emb_ckmux2m8(A, B, S, Z);
input  A;
input  B;
input  S;
output Z;

assign Z = S ? B : A;

endmodule

module gclk_clk_gate(
                 gate_en ,
                 clk_gate_in ,
                 test_mode ,
                 clk_gate_out
);
input            gate_en ;
input            clk_gate_in ;
input            test_mode ;

output           clk_gate_out;

reg q;
always @ (*) begin
    if (clk_gate_in==1'b0)
     q = test_mode||gate_en ;
end
assign clk_gate_out = clk_gate_in & q;

endmodule

//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_clkgate(
                      test_mode    ,
                      clk          ,
                      ce_pra       ,
                      ce_mult_u    ,
                      ce_mult_l    ,
                      ce_poa       ,
                      ce_comp      ,
                      ce_ufc       ,
                      ce_ibuf      ,
                      clk_pra      ,
                      clk_mult_u   ,
                      clk_mult_l   ,
                      clk_poa      ,
                      clk_comp     ,
                      clk_ufc      ,
                      clk_ibuf      
                  );
input   test_mode    ;
input   clk          ;
input   ce_pra       ;
input   ce_mult_u    ;
input   ce_mult_l    ;
input   ce_poa       ;
input   ce_comp      ;
input   ce_ufc       ;
input   ce_ibuf      ;

output  clk_pra      ;
output  clk_mult_u   ;
output  clk_mult_l   ;
output  clk_poa      ;
output  clk_comp     ;
output  clk_ufc      ;
output  clk_ibuf     ;


gclk_clk_gate U_gclk_clk_gate_pra (
                .test_mode       (test_mode  ),       
                .clk_gate_in     (clk        ),         
                .gate_en         (ce_pra     ),     
                .clk_gate_out    (clk_pra    )      
);


//----------------------------------------------
gclk_clk_gate U_gclk_clk_gate_mult_u (
                .test_mode       (test_mode     ),       
                .clk_gate_in     (clk           ),         
                .gate_en         (ce_mult_u     ),     
                .clk_gate_out    (clk_mult_u    )      
);



//----------------------------------------------
gclk_clk_gate U_gclk_clk_gate_mult_l (
                .test_mode       (test_mode     ),       
                .clk_gate_in     (clk           ),         
                .gate_en         (ce_mult_l     ),     
                .clk_gate_out    (clk_mult_l    )      
);


//----------------------------------------------
gclk_clk_gate U_gclk_clk_gate_poa (
                .test_mode       (test_mode     ),       
                .clk_gate_in     (clk           ),         
                .gate_en         (ce_poa     ),     
                .clk_gate_out    (clk_poa    )      
);


//----------------------------------------------
gclk_clk_gate U_gclk_clk_gate_comp (
                .test_mode       (test_mode     ),       
                .clk_gate_in     (clk           ),         
                .gate_en         (ce_comp     ),     
                .clk_gate_out    (clk_comp    )      
);


//----------------------------------------------
gclk_clk_gate U_gclk_clk_gate_ufc (
                .test_mode       (test_mode     ),       
                .clk_gate_in     (clk           ),         
                .gate_en         (ce_ufc     ),     
                .clk_gate_out    (clk_ufc    )      
);


//----------------------------------------------
gclk_clk_gate U_gclk_clk_gate_ibuf (
                .test_mode       (test_mode     ),       
                .clk_gate_in     (clk           ),         
                .gate_en         (ce_ibuf     ),     
                .clk_gate_out    (clk_ibuf    )      
);

endmodule
//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_compunit(
                       clk_comp        ,                          
                       rst_n      ,                            
                       R_pre      ,                            
                       U_buf      ,                            
                       cfg_vldbit ,                                 
                       cfg_match  ,                                
                       cfg_imatch ,                                 
                       MATCH      ,                            
                       UNDERFLOW  ,                                
                       iMATCH     ,    
                       OVERFLOW        
                                          );

//clock and reset
input           clk_comp;
input           rst_n;   //sys reset

input  [55:0]   R_pre;  
input  [55:0]   U_buf;  
input  [55:0]   cfg_vldbit;
input           cfg_match;
input           cfg_imatch;

output          MATCH;
output          UNDERFLOW;
output          iMATCH;
output          OVERFLOW;
wire   [55:0]   w56_comp_r;
wire   [55:0]   w56_comp_u;
wire   [55:0]   w56_comp_ub;

reg             match_0;
reg             match_1;
reg             imatch_0;
reg             imatch_1;

DSPCELL_AND2 #(56) U_DSPCELL_AND2_COMP_R ( //assign o = i0 & i1;
                        .i0  (cfg_vldbit  ),
                        .i1  (R_pre       ),
                        .o   (w56_comp_r  ) 
);
DSPCELL_AND2 #(56) U_DSPCELL_AND2_COMP_U ( //assign o = i0 & i1;
                        .i0  (cfg_vldbit  ),
                        .i1  (U_buf       ),
                        .o   (w56_comp_u  ) 
);
DSPCELL_AND2 #(56) U_DSPCELL_AND2_COMP_UB ( //assign o = i0 & i1;
                        .i0  (cfg_vldbit  ),
                        .i1  (~U_buf       ),
                        .o   (w56_comp_ub  ) 
);
always @(posedge clk_comp or negedge rst_n) begin
   if(rst_n == 0) begin
       match_0 <= `DLY 0;
   end
   else if(w56_comp_r == w56_comp_u) begin
       match_0 <= `DLY 1;
   end
   else begin
       match_0 <= `DLY 0;
   end
end
always @(posedge clk_comp or negedge rst_n) begin
   if(rst_n == 0) begin
       imatch_0 <= `DLY 0;
   end
   else if(w56_comp_r == w56_comp_ub) begin
       imatch_0 <= `DLY 1;
   end
   else begin
       imatch_0 <= `DLY 0;
   end
end
always @(posedge clk_comp or negedge rst_n) begin
   if(rst_n == 0) begin
       match_1  <= `DLY 0;
       imatch_1 <= `DLY 0;
   end
   else begin
       match_1  <= `DLY match_0 ;
       imatch_1 <= `DLY imatch_0;
   end
end
DSPCELL_MUX2 #(1) U_DSPCELL_MUX2_COMP_M(
                .i0   (match_1     ),
                .i1   (match_0     ),
                .sel  (cfg_match   ),
                .o    (MATCH       )
);
DSPCELL_MUX2 #(1) U_DSPCELL_MUX2_COMP_iM(
                .i0   (imatch_1     ),
                .i1   (imatch_0     ),
                .sel  (cfg_imatch   ),
                .o    (iMATCH       )
);

DSPCELL_AND3 #(1) U_DSPCELL_AND3_COMP_UDFL (
                .i0 (~match_0   ),
                .i1 (~imatch_0  ),
                .i2 (match_1    ),
                .o  (UNDERFLOW  ) 
);

DSPCELL_AND3 #(1) U_DSPCELL_AND3_COMP_OVFL (
                .i0 (~match_0   ),
                .i1 (~imatch_0  ),
                .i2 (imatch_1   ),
                .o  (OVERFLOW   ) 
);

endmodule

// VPERL: GENERATED_BEG

module dsp_core (
	alcasout,
	aucasout,
	clcasout,
	cucasout,
	imatch,
	match,
	overflow,
	r,
	rcarrycasout,
	rcasout,
	recarrycasout,
	underflow,
	al,
	alcasin,
	au,
	aucasin,
	cecomp,
	ceibuf,
	cemultl,
	cemultu,
	cepoa,
	cepra,
	ceufc,
	cfg_aluctrl,
	cfg_blctrl,
	cfg_buctrl,
	cfg_cctrl,
	cfg_fcctrl,
	cfg_frctrl,
	cfg_imatch,
	cfg_mat_clr,
	cfg_match,
	cfg_mctrl,
	cfg_mult_l,
	cfg_mult_u,
	cfg_parctrl,
	cfg_pasctrl,
	cfg_pasubctrl,
	cfg_pazctrl,
	cfg_poa_ceyin,
	cfg_poa_ceyout,
	cfg_poa_cyout,
	cfg_poa_rout,
	cfg_pra_al,
	cfg_pra_au,
	cfg_pra_cl,
	cfg_pra_cu,
	cfg_pra_dl,
	cfg_pra_du,
	cfg_pra_ol,
	cfg_pra_ou,
	cfg_rndm,
	cfg_subctrl,
	cfg_ufcctrl,
	cfg_ufcmux,
	cfg_vldbit,
	cl,
	clcasin,
	clk,
	cu,
	cucasin,
	dl,
	du,
	ialuctrl,
	iblctrl,
	ibuctrl,
	icctrl,
	ifcctrl,
	ifrctrl,
	imctrl,
	iparctrl,
	ipasctrl,
	ipasubctrl,
	ipazctrl,
	irndm,
	isubctrl,
	iufcctrl,
	rcarrycasin,
	rcasin,
	recarrycasin,
	rstn,
	sck,
	sen,
	si,
	smode,
	srst,
	u 
);

output	[17:0]	alcasout;
output	[17:0]	aucasout;
output	[17:0]	clcasout;
output	[17:0]	cucasout;
output		imatch;
output		match;
output		overflow;
output	[71:0]	r;
output		rcarrycasout;
output	[55:0]	rcasout;
output		recarrycasout;
output		underflow;
input	[17:0]	al;
input	[17:0]	alcasin;
input	[17:0]	au;
input	[17:0]	aucasin;
input		cecomp;
input		ceibuf;
input		cemultl;
input		cemultu;
input		cepoa;
input		cepra;
input		ceufc;
input		cfg_aluctrl;
input		cfg_blctrl;
input		cfg_buctrl;
input		cfg_cctrl;
input		cfg_fcctrl;
input		cfg_frctrl;
input		cfg_imatch;
input		cfg_mat_clr;
input		cfg_match;
input		cfg_mctrl;
input	[1:0]	cfg_mult_l;
input	[1:0]	cfg_mult_u;
input		cfg_parctrl;
input		cfg_pasctrl;
input		cfg_pasubctrl;
input		cfg_pazctrl;
input		cfg_poa_ceyin;
input		cfg_poa_ceyout;
input		cfg_poa_cyout;
input	[1:0]	cfg_poa_rout;
input	[2:0]	cfg_pra_al;
input	[2:0]	cfg_pra_au;
input	[2:0]	cfg_pra_cl;
input	[2:0]	cfg_pra_cu;
input		cfg_pra_dl;
input		cfg_pra_du;
input		cfg_pra_ol;
input		cfg_pra_ou;
input		cfg_rndm;
input		cfg_subctrl;
input		cfg_ufcctrl;
input		cfg_ufcmux;
input	[55:0]	cfg_vldbit;
input	[17:0]	cl;
input	[17:0]	clcasin;
input		clk;
input	[17:0]	cu;
input	[17:0]	cucasin;
input	[17:0]	dl;
input	[17:0]	du;
input	[2:0]	ialuctrl;
input		iblctrl;
input		ibuctrl;
input	[2:0]	icctrl;
input	[2:0]	ifcctrl;
input	[1:0]	ifrctrl;
input	[5:0]	imctrl;
input	[5:0]	iparctrl;
input	[7:0]	ipasctrl;
input	[1:0]	ipasubctrl;
input	[5:0]	ipazctrl;
input		irndm;
input	[2:0]	isubctrl;
input		iufcctrl;
input		rcarrycasin;
input	[55:0]	rcasin;
input		recarrycasin;
input		rstn;
input		sck;
input		sen;
input		si;
input		smode;
input		srst;
input	[55:0]	u;

wire	[2:0]	aluctrl;
wire		blctrl;
wire		buctrl;
wire	[2:0]	cctrl;
wire		clk_comp;
wire		clk_ibuf;
wire		clk_mult_l;
wire		clk_mult_u;
wire		clk_poa;
wire		clk_pra;
wire		clk_ufc;
wire	[2:0]	fcctrl;
wire	[1:0]	frctrl;
wire	[17:0]	mal;
wire	[17:0]	mau;
wire	[17:0]	mbl;
wire	[17:0]	mbu;
wire	[5:0]	mctrl;
wire	[55:0]	mrl;
wire	[55:0]	mru;
wire	[5:0]	parctrl;
wire	[7:0]	pasctrl;
wire	[1:0]	pasubctrl;
wire	[5:0]	pazctrl;
wire		rndm;
wire	[55:0]	rpre;
wire	[2:0]	subctrl;
wire	[55:0]	ubuf;
wire	[55:0]	ufc;
wire		ufcctrl;

dsp_clkgate U_dsp_clkgate (
	.test_mode	(smode),
	.clk		(clk),
	.ce_pra		(cepra),
	.ce_mult_u	(cemultu),
	.ce_mult_l	(cemultl),
	.ce_poa		(cepoa),
	.ce_comp	(cecomp),
	.ce_ufc		(ceufc),
	.ce_ibuf	(ceibuf),

	.clk_pra	(clk_pra),
	.clk_mult_u	(clk_mult_u),
	.clk_mult_l	(clk_mult_l),
	.clk_poa	(clk_poa),
	.clk_comp	(clk_comp),
	.clk_ufc	(clk_ufc),
	.clk_ibuf	(clk_ibuf) 
);

dsp_compunit U_dsp_compunit (
	.clk_comp	(clk_comp),
	.rst_n		(rstn),
	.R_pre		(rpre[55:0]),
	.U_buf		(ubuf[55:0]),
	.cfg_vldbit	(cfg_vldbit[55:0]),
	.cfg_match	(cfg_match),
	.cfg_imatch	(cfg_imatch),

	.MATCH		(match),
	.UNDERFLOW	(underflow),
	.iMATCH		(imatch),
	.OVERFLOW	(overflow) 
);

dsp_input_buf U_dsp_input_buf (
	.clk_ibuf	(clk_ibuf),
	.rst_n		(rstn),
	.cfg_PAZCTRL	(cfg_pazctrl),
	.cfg_PARCTRL	(cfg_parctrl),
	.cfg_PASUBCTRL	(cfg_pasubctrl),
	.cfg_BLCTRL	(cfg_blctrl),
	.cfg_BUCTRL	(cfg_buctrl),
	.cfg_PASCTRL	(cfg_pasctrl),
	.cfg_ALUCTRL	(cfg_aluctrl),
	.cfg_FCCTRL	(cfg_fcctrl),
	.cfg_UFCCTRL	(cfg_ufcctrl),
	.cfg_SUBCTRL	(cfg_subctrl),
	.cfg_MCTRL	(cfg_mctrl),
	.cfg_CCTRL	(cfg_cctrl),
	.cfg_FRCTRL	(cfg_frctrl),
	.cfg_RNDM	(cfg_rndm),
	.iPAZCTRL	(ipazctrl[5:0]),
	.iPARCTRL	(iparctrl[5:0]),
	.iPASUBCTRL	(ipasubctrl[1:0]),
	.iBLCTRL	(iblctrl),
	.iBUCTRL	(ibuctrl),
	.iPASCTRL	(ipasctrl[7:0]),
	.iALUCTRL	(ialuctrl[2:0]),
	.iFCCTRL	(ifcctrl[2:0]),
	.iUFCCTRL	(iufcctrl),
	.iSUBCTRL	(isubctrl[2:0]),
	.iMCTRL		(imctrl[5:0]),
	.iCCTRL		(icctrl[2:0]),
	.iFRCTRL	(ifrctrl[1:0]),
	.iRNDM		(irndm),

	.PAZCTRL	(pazctrl[5:0]),
	.PARCTRL	(parctrl[5:0]),
	.PASUBCTRL	(pasubctrl[1:0]),
	.BLCTRL		(blctrl),
	.BUCTRL		(buctrl),
	.PASCTRL	(pasctrl[7:0]),
	.ALUCTRL	(aluctrl[2:0]),
	.FCCTRL		(fcctrl[2:0]),
	.UFCCTRL	(ufcctrl),
	.SUBCTRL	(subctrl[2:0]),
	.MCTRL		(mctrl[5:0]),
	.CCTRL		(cctrl[2:0]),
	.FRCTRL		(frctrl[1:0]),
	.RNDM		(rndm) 
);

dsp_multblock U_dsp_multblock (
	.clk_mult_u	(clk_mult_u),
	.clk_mult_l	(clk_mult_l),
	.rst_n		(rstn),
	.MA_U		(mau[17:0]),
	.MB_U		(mbu[17:0]),
	.MA_L		(mal[17:0]),
	.MB_L		(mbl[17:0]),
	.U_buf		(ubuf[55:0]),
	.R		(r[55:0]),
	.cfg_mult_u	(cfg_mult_u[1:0]),
	.cfg_mult_l	(cfg_mult_l[1:0]),
	.MCTRL		(mctrl[5:0]),

	.MR_U		(mru[55:0]),
	.MR_L		(mrl[55:0]) 
);

dsp_postadder U_dsp_postadder (
	.clk_poa		(clk_poa),
	.rst_n			(rstn),
	.MR_U			(mru[55:0]),
	.MR_L			(mrl[55:0]),
	.UFC			(ufc[55:0]),
	.R_CARRY_CAS_IN		(rcarrycasin),
	.R_ECARRY_CAS_IN	(recarrycasin),
	.MATCH			(match),
	.RNDM			(rndm),
	.SUBCTRL		(subctrl[2:0]),
	.ALUCTRL		(aluctrl[2:0]),
	.FRCTRL			(frctrl[1:0]),
	.CCTRL			(cctrl[2:0]),
	.cfg_mat_clr		(cfg_mat_clr),
	.cfg_poa_cyout		(cfg_poa_cyout),
	.cfg_poa_ceyout		(cfg_poa_ceyout),
	.cfg_poa_ceyin		(cfg_poa_ceyin),
	.cfg_poa_rout		(cfg_poa_rout[1:0]),

	.R_CARRY_CAS_OUT	(rcarrycasout),
	.R_ECARRY_CAS_OUT	(recarrycasout),
	.R_pre			(rpre[55:0]),
	.R			(r[71:0]),
	.R_CAS_OUT		(rcasout[55:0]) 
);

dsp_preadder U_dsp_preadder (
	.clk_pra	(clk_pra),
	.rst_n		(rstn),
	.A_L		(al[17:0]),
	.C_L		(cl[17:0]),
	.D_L		(dl[17:0]),
	.A_U		(au[17:0]),
	.C_U		(cu[17:0]),
	.D_U		(du[17:0]),
	.A_L_CAS_IN	(alcasin[17:0]),
	.C_L_CAS_IN	(clcasin[17:0]),
	.A_U_CAS_IN	(aucasin[17:0]),
	.C_U_CAS_IN	(cucasin[17:0]),
	.PAZCTRL	(pazctrl[5:0]),
	.PARCTRL	(parctrl[5:0]),
	.PASUBCTRL	(pasubctrl[1:0]),
	.BLCTRL		(blctrl),
	.BUCTRL		(buctrl),
	.PASCTRL	(pasctrl[7:0]),
	.cfg_pra_au	(cfg_pra_au[2:0]),
	.cfg_pra_cu	(cfg_pra_cu[2:0]),
	.cfg_pra_du	(cfg_pra_du),
	.cfg_pra_dl	(cfg_pra_dl),
	.cfg_pra_al	(cfg_pra_al[2:0]),
	.cfg_pra_cl	(cfg_pra_cl[2:0]),
	.cfg_pra_ou	(cfg_pra_ou),
	.cfg_pra_ol	(cfg_pra_ol),

	.A_L_CAS_OUT	(alcasout[17:0]),
	.C_L_CAS_OUT	(clcasout[17:0]),
	.A_U_CAS_OUT	(aucasout[17:0]),
	.C_U_CAS_OUT	(cucasout[17:0]),
	.MA_U		(mau[17:0]),
	.MB_U		(mbu[17:0]),
	.MB_L		(mbl[17:0]),
	.MA_L		(mal[17:0]) 
);

dsp_ufcmux U_dsp_ufcmux (
	.clk_ufc	(clk_ufc),
	.rst_n		(rstn),
	.R_CAS_IN	(rcasin[55:0]),
	.R		(r[55:0]),
	.U		(u[55:0]),
	.FCCTRL		(fcctrl[2:0]),
	.UFCCTRL	(ufcctrl),
	.cfg_ufcmux	(cfg_ufcmux),

	.UFC		(ufc[55:0]),
	.U_BUF		(ubuf[55:0]) 
);

endmodule

// VPERL: GENERATED_END

//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_input_buf(
                clk_ibuf,
                rst_n,   //sys reset
                cfg_PAZCTRL   ,    //             
                cfg_PARCTRL   ,    //             
                cfg_PASUBCTRL ,    //               
                cfg_BLCTRL    ,    //            
                cfg_BUCTRL    ,    //            
                cfg_PASCTRL   ,    //             
                cfg_ALUCTRL   ,    //   I Input Control the functionality of ALU operation 
                cfg_FCCTRL    ,    //   I Input Select Feedback and Cascaded data for UFC MUX 
                cfg_UFCCTRL   ,    //   I Input Select U and FC MUX data for post stage operation
                cfg_SUBCTRL   ,    //   I Input Select and Control to perform Subtraction in post stage operation 
                cfg_MCTRL     ,    //   I Input Select and Control the result of lower and upper multipliers and source for MR_U MUX 
                cfg_CCTRL     ,    //   I Input Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
                cfg_FRCTRL    ,    //   I Input Select final result source 
                cfg_RNDM      ,    //   I Input Rounding method from user logic: 0 Rounding to Zero, 1:Rounding to infinity 
                iPAZCTRL   ,    //             
                iPARCTRL   ,    //             
                iPASUBCTRL ,    //               
                iBLCTRL    ,    //            
                iBUCTRL    ,    //            
                iPASCTRL   ,    //             
                iALUCTRL   ,    //   I Input Control the functionality of ALU operation 
                iFCCTRL    ,    //   I Input Select Feedback and Cascaded data for UFC MUX 
                iUFCCTRL   ,    //   I Input Select U and FC MUX data for post stage operation
                iSUBCTRL   ,    //   I Input Select and Control to perform Subtraction in post stage operation 
                iMCTRL     ,    //   I Input Select and Control the result of lower and upper multipliers and source for MR_U MUX 
                iCCTRL     ,    //   I Input Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
                iFRCTRL    ,    //   I Input Select final result source 
                iRNDM      ,    //   I Input Rounding method from user logic: 0 Rounding to Zero, 1:Rounding to infinity 
                
                PAZCTRL   ,    //             
                PARCTRL   ,    //             
                PASUBCTRL ,    //               
                BLCTRL    ,    //            
                BUCTRL    ,    //            
                PASCTRL   ,    //             
                ALUCTRL   ,    //   I Input Control the functionality of ALU operation 
                FCCTRL    ,    //   I Input Select Feedback and Cascaded data for UFC MUX 
                UFCCTRL   ,    //   I Input Select U and FC MUX data for post stage operation
                SUBCTRL   ,    //   I Input Select and Control to perform Subtraction in post stage operation 
                MCTRL     ,    //   I Input Select and Control the result of lower and upper multipliers and source for MR_U MUX 
                CCTRL     ,    //   I Input Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
                FRCTRL    ,    //   I Input Select final result source 
                RNDM           //   I Input Rounding method from user logic: 0 Rounding to Zero, 1:Rounding to infinity 



                     
                  );

 

//clock and reset
input              clk_ibuf;
input              rst_n;   //sys reset
                            //iPACTRL   24  I Input Select and Control the functionality of the Pre-Adder and Selector
input              cfg_PAZCTRL   ;    //             
input              cfg_PARCTRL   ;    //             
input              cfg_PASUBCTRL ;    //               
input              cfg_BLCTRL    ;    //            
input              cfg_BUCTRL    ;    //            
input              cfg_PASCTRL   ;    //             
input              cfg_ALUCTRL   ;    //   I Input Control the functionality of ALU operation 
input              cfg_FCCTRL    ;    //   I Input Select Feedback and Cascaded data for UFC MUX 
input              cfg_UFCCTRL   ;    //   I Input Select U and FC MUX data for post stage operation
input              cfg_SUBCTRL   ;    //   I Input Select and Control to perform Subtraction in post stage operation 
input              cfg_MCTRL     ;    //   I Input Select and Control the result of lower and upper multipliers and source for MR_U MUX 
input              cfg_CCTRL     ;    //   I Input Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
input              cfg_FRCTRL    ;    //   I Input Select final result source 
input              cfg_RNDM      ;    //   I Input Rounding method from user logic: 0 Rounding to Zero, 1:Rounding to infinity 

input      [5:0 ]  iPAZCTRL   ;    //             
input      [5:0 ]  iPARCTRL   ;    //             
input      [1:0 ]  iPASUBCTRL ;    //               
input              iBLCTRL    ;    //            
input              iBUCTRL    ;    //            
input      [7:0 ]  iPASCTRL   ;    //             
input      [2:0 ]  iALUCTRL   ;    //   I Input Control the functionality of ALU operation 
input      [2:0 ]  iFCCTRL    ;    //   I Input Select Feedback and Cascaded data for UFC MUX 
input              iUFCCTRL   ;    //   I Input Select U and FC MUX data for post stage operation
input      [2:0 ]  iSUBCTRL   ;    //   I Input Select and Control to perform Subtraction in post stage operation 
input      [5:0 ]  iMCTRL     ;    //   I Input Select and Control the result of lower and upper multipliers and source for MR_U MUX 
input      [2:0 ]  iCCTRL     ;    //   I Input Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
input      [1:0 ]  iFRCTRL    ;    //   I Input Select final result source 
input              iRNDM      ;    //   I Input Rounding method from user logic: 0 Rounding to Zero, 1:Rounding to infinity 

output     [5:0 ]  PAZCTRL   ;    //             
output     [5:0 ]  PARCTRL   ;    //             
output     [1:0 ]  PASUBCTRL ;    //               
output             BLCTRL    ;    //            
output             BUCTRL    ;    //            
output     [7:0 ]  PASCTRL   ;    //             
output     [2:0 ]  ALUCTRL   ;    //   I Input Control the functionality of ALU operation 
output     [2:0 ]  FCCTRL    ;    //   I Input Select Feedback and Cascaded data for UFC MUX 
output             UFCCTRL   ;    //   I Input Select U and FC MUX data for post stage operation
output     [2:0 ]  SUBCTRL   ;    //   I Input Select and Control to perform Subtraction in post stage operation 
output     [5:0 ]  MCTRL     ;    //   I Input Select and Control the result of lower and upper multipliers and source for MR_U MUX 
output     [2:0 ]  CCTRL     ;    //   I Input Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
output     [1:0 ]  FRCTRL    ;    //   I Input Select final result source 
output             RNDM      ;    //   I Input Rounding method from user logic: 0 Rounding to Zero, 1:Rounding to infinity 




DSPCELL_SELBUF #(6)  U_DSPCELL_SELBUF_IBUF0 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iPAZCTRL         ),
                     .sel      (cfg_PAZCTRL      ),
                     .o        (PAZCTRL          ) 
);
DSPCELL_SELBUF #(6)  U_DSPCELL_SELBUF_IBUF1 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iPARCTRL         ),
                     .sel      (cfg_PARCTRL      ),
                     .o        (PARCTRL          ) 
);

DSPCELL_SELBUF #(2)  U_DSPCELL_SELBUF_IBUF2 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iPASUBCTRL         ),
                     .sel      (cfg_PASUBCTRL      ),
                     .o        (PASUBCTRL          ) 
);
DSPCELL_SELBUF #(1)  U_DSPCELL_SELBUF_IBUF3 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iBLCTRL         ),
                     .sel      (cfg_BLCTRL      ),
                     .o        (BLCTRL          ) 
);
DSPCELL_SELBUF #(1)  U_DSPCELL_SELBUF_IBUF4 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iBUCTRL         ),
                     .sel      (cfg_BUCTRL      ),
                     .o        (BUCTRL          ) 
);
DSPCELL_SELBUF #(8)  U_DSPCELL_SELBUF_IBUF5 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iPASCTRL         ),
                     .sel      (cfg_PASCTRL      ),
                     .o        (PASCTRL          ) 
);
DSPCELL_SELBUF #(3)  U_DSPCELL_SELBUF_IBUF6 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iALUCTRL         ),
                     .sel      (cfg_ALUCTRL      ),
                     .o        (ALUCTRL          ) 
);
DSPCELL_SELBUF #(3)  U_DSPCELL_SELBUF_IBUF7 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iFCCTRL         ),
                     .sel      (cfg_FCCTRL      ),
                     .o        (FCCTRL          ) 
);
DSPCELL_SELBUF #(1)  U_DSPCELL_SELBUF_IBUF8 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iUFCCTRL         ),
                     .sel      (cfg_UFCCTRL      ),
                     .o        (UFCCTRL          ) 
);
DSPCELL_SELBUF #(3)  U_DSPCELL_SELBUF_IBUF9 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iSUBCTRL         ),
                     .sel      (cfg_SUBCTRL      ),
                     .o        (SUBCTRL          ) 
);
DSPCELL_SELBUF #(6)  U_DSPCELL_SELBUF_IBUF10 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iMCTRL         ),
                     .sel      (cfg_MCTRL      ),
                     .o        (MCTRL          ) 
);
DSPCELL_SELBUF #(3)  U_DSPCELL_SELBUF_IBUF11 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iCCTRL         ),
                     .sel      (cfg_CCTRL      ),
                     .o        (CCTRL          ) 
);
DSPCELL_SELBUF #(2)  U_DSPCELL_SELBUF_IBUF12 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iFRCTRL         ),
                     .sel      (cfg_FRCTRL      ),
                     .o        (FRCTRL          ) 
);
DSPCELL_SELBUF #(1)  U_DSPCELL_SELBUF_IBUF13 (  
                     .clk      (clk_ibuf              ),
                     .rst_n    (rst_n            ),  
                     .i        (iRNDM         ),
                     .sel      (cfg_RNDM      ),
                     .o        (RNDM          ) 
);


endmodule
//*************************************************
//author:    hywang
//date:      20140522
//function:   1)DSPCELL common cell
//            2)
//*************************************************
//$Log: .v,v $

`ifdef DLY_DSP
`else
`define DLY_DSP #0.1
`endif

`ifdef DLY
`else
`define DLY #0.1
`endif




//==========================================================
module DSPCELL_AND2 ( //assign o = i0 & i1;
      i0,
      i1,
      o  
);
parameter WIDTH = 1;
input [WIDTH-1:0]  i0;
input [WIDTH-1:0]  i1;
output[WIDTH-1:0]  o;

`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
	assign o = i0 & i1;
`endif
endmodule
//==========================================================

module DSPCELL_AND3 (
    i0,
    i1,
    i2,
    o  
);
parameter WIDTH = 1;
input  [WIDTH-1:0] i0;
input  [WIDTH-1:0] i1;
input  [WIDTH-1:0] i2;
output [WIDTH-1:0] o;
`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
	assign o = i0 & i1 & i2;
`endif
endmodule
//==========================================================
module DSPCELL_MUX2(  //assign o = sel ? i1 : i0;
                      i0,        
                      i1,     
                      sel,    
                      o         
);
parameter WIDTH = 1;
input [WIDTH-1:0] i0;
input [WIDTH-1:0] i1;
input             sel;
output[WIDTH-1:0] o;


`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
	assign o = sel ? i1 : i0;
//genvar i; 
//generate for(i=0; i<WIDTH; i=i+1) begin:gmux2
//gclk_clk_mux U_gclk_clk_mux(
//      .ck_i0      (i0[i]  ),
//      .ck_i1      (i1[i]  ),
//      .sel        (sel     ),
//      .ck_out     (o[i] )
//);
//end
//endgenerate
`endif
endmodule
//==========================================================
//==========================================================
module DSPCELL_MUX4(  
                      i0,        
                      i1,     
                      i2,     
                      i3,     
                      sel,    
                      o         
);
parameter WIDTH = 1;
input [WIDTH-1:0] i0;
input [WIDTH-1:0] i1;
input [WIDTH-1:0] i2;
input [WIDTH-1:0] i3;
input [1:0]       sel;
output[WIDTH-1:0] o;

wire  [WIDTH-1:0] o_0;
wire  [WIDTH-1:0] o_1;

`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
DSPCELL_MUX2 #(WIDTH) U_DSPCELL_MUX2_0(
                .i0   (i0     ),  
                .i1   (i1     ),  
                .sel  (sel[0] ),   
                .o    (o_0    )  
);
DSPCELL_MUX2 #(WIDTH) U_DSPCELL_MUX2_1(
                .i0   (i2     ),  
                .i1   (i3     ),  
                .sel  (sel[0] ),   
                .o    (o_1    )  
);
DSPCELL_MUX2 #(WIDTH) U_DSPCELL_MUX2_2(
                .i0   (o_0     ),  
                .i1   (o_1     ),  
                .sel  (sel[1]  ),   
                .o    (o       )  
);

`endif
endmodule
//==========================================================
module DSPCELL_MUX8(  
                      i0,        
                      i1,     
                      i2,     
                      i3,     
                      i4,     
                      i5,     
                      i6,     
                      i7,     
                      sel,    
                      o         
);
parameter WIDTH = 1;
input [WIDTH-1:0] i0;
input [WIDTH-1:0] i1;
input [WIDTH-1:0] i2;
input [WIDTH-1:0] i3;
input [WIDTH-1:0] i4;
input [WIDTH-1:0] i5;
input [WIDTH-1:0] i6;
input [WIDTH-1:0] i7;
input [2:0]       sel;
output[WIDTH-1:0] o;

wire  [WIDTH-1:0] o_0;
wire  [WIDTH-1:0] o_1;

`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
DSPCELL_MUX4 #(WIDTH) U_DSPCELL_MUX4_0(
                .i0   (i0     ),  
                .i1   (i1     ),  
                .i2   (i2     ),  
                .i3   (i3     ),  
                .sel  (sel[1:0] ),   
                .o    (o_0    )  
);
DSPCELL_MUX4 #(WIDTH) U_DSPCELL_MUX4_1(
                .i0   (i4     ),  
                .i1   (i5     ),  
                .i2   (i6     ),  
                .i3   (i7     ),  
                .sel  (sel[1:0] ),   
                .o    (o_1    )  
);
DSPCELL_MUX2 #(WIDTH) U_DSPCELL_MUX2_2(
                .i0   (o_0     ),  
                .i1   (o_1     ),  
                .sel  (sel[2]  ),   
                .o    (o       )  
);

`endif
endmodule
//==========================================================



module DSPCELL_SELBUF(  //assign o = sel == 0 ? o_buf :  i
                      clk,        
                      rst_n,
                      i,     
                      sel,    
                      o         
);
parameter WIDTH = 1;
input             clk;
input             rst_n;
input [WIDTH-1:0] i;
input             sel;
output[WIDTH-1:0] o;
reg   [WIDTH-1:0] o_buf;
`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
always @(posedge clk or negedge rst_n) begin
    if(rst_n == 0) begin
        o_buf <= 0;
    end
    else begin
        o_buf <= i;
    end
end
assign o = sel == 0 ? o_buf :  i;
`endif

endmodule
//==========================================================
module DSPCELL_FULLADD(  //s = i0 + i1
                      i0,        
                      i1,     
                      s,    
                      ci,         
                      co         
);
parameter WIDTH = 1;
input [WIDTH-1:0] i0;
input [WIDTH-1:0] i1;
input             ci;
output[WIDTH-1:0] s;
output            co;
wire  [WIDTH:0]   s_temp;
`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
assign  `DLY_DSP s_temp = i0 + i1 + ci;
assign s = s_temp[WIDTH-1:0];
assign co = s_temp[WIDTH];
`endif

endmodule

//==========================================================
module DSPCELL_ADD(  //s = i0 + i1
                      i0,        
                      i1,     
                      s,    
                      c         
);
parameter WIDTH = 1;
input [WIDTH-1:0] i0;
input [WIDTH-1:0] i1;
output[WIDTH-1:0] s;
output            c;
wire  [WIDTH:0]   s_temp;
`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
assign  `DLY_DSP s_temp = i0 + i1;
assign s = s_temp[WIDTH-1:0];
assign c = s_temp[WIDTH];
`endif

endmodule
//==========================================================
module DSPCELL_BIT_ADD(  
                      i0,        
                      i1,     
                      i2,     
                      s,
                      c    
);
parameter WIDTH = 1;

input   [WIDTH-1:0]   i0;
input   [WIDTH-1:0]   i1;
input   [WIDTH-1:0]   i2;
output  [WIDTH-1:0]   s;
output  [WIDTH-1:0]   c;
wire    [WIDTH*2-1:0] temp;
`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
generate
genvar i;
for(i =0;i<WIDTH;i = i + 1) 
begin: adder
   assign temp[i*2+1:i*2] = i0[i] + i1[i] + i2[i];
   assign `DLY_DSP s[i] = temp[i*2];
   assign `DLY_DSP c[i] = temp[i*2+1];
end
endgenerate
`endif
endmodule


/*
//==========================================================
module DSPCELL_SUB(  // s = i0 - i1 
                      i0,        
                      i1,     
                      s,    
                      c         
);
parameter WIDTH = 1;
input [WIDTH-1:0] i0;
input [WIDTH-1:0] i1;
output[WIDTH-1:0] s;
output            c;
wire  [WIDTH:0]   s_temp;
`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
assign s_temp = i0 - i1;
assign `DLY_DSP s = s_temp[WIDTH-1:0];
assign `DLY_DSP c = s_temp[WIDTH];
`endif
endmodule
*/
//==========================================================
module DSPCELL_MULT(  // s = i0 * i1 
                      i0,        
                      i1,     
                      o    
);
parameter WIDTH = 1;

input   [WIDTH-1:0]   i0;
input   [WIDTH-1:0]   i1;
output  [WIDTH*2-1:0] o;
wire signed  [WIDTH-1:0]    i0;
wire signed  [WIDTH-1:0]    i1;
wire signed  [WIDTH*2-1:0]  o;

`ifdef   DSPCELL_GATE
   `ifdef UMC55SP
   `elsif UMC40LP
   `endif
`else
assign `DLY_DSP o = i0 * i1;
`endif
endmodule
//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_multblock(
                         clk_mult_u, 
                         clk_mult_l, 
                         rst_n,
                         MA_U ,   
                         MB_U ,   
                         MA_L ,   
                         MB_L ,   
                         U_buf,  
                         R,  
                         MR_U ,   
                         MR_L ,     
                         cfg_mult_u,
                         cfg_mult_l,
                         MCTRL         
                                     );

 

//clock and reset
input           clk_mult_u;
input           clk_mult_l;
input           rst_n;   //sys reset

input  [17:0]   MA_U;  
input  [17:0]   MB_U;  
input  [17:0]   MA_L;  
input  [17:0]   MB_L;  
input  [55:0]   U_buf;  
input  [55:0]   R;  

output [55:0]   MR_U;  
output [55:0]   MR_L;  

input  [1:0]    cfg_mult_u;
input  [1:0]    cfg_mult_l;
input  [5:0]    MCTRL;

wire   [35:0]   w36_mabu;
wire   [35:0]   w36_mabu1;
wire   [35:0]   w36_mabu2;
wire   [35:0]   w36_mabu3;
wire   [52:0]   w53_mabu4;

wire   [35:0]   w36_mabl;
wire   [35:0]   w36_mabl1;
wire   [35:0]   w36_mabl2;
wire   [35:0]   w36_mabl3;

wire   [55:0]   w56_mcat;
wire   [55:0]   MR_L_t;

DSPCELL_MULT #(18) U_DSPCELL_MULT_MABU0(
                     .i0 (MA_U      ),
                     .i1 (MB_U      ),
                     .o  (w36_mabu  ) 
);
DSPCELL_SELBUF #(36) U_DSPCELL_SELBUF_U1(  //assign o = sel == 0 ? o_buf :  i
                     .clk  (clk_mult_u           ),       
                     .rst_n(rst_n         ),       
                     .i    (w36_mabu      ),     
                     .sel  (cfg_mult_u[0] ),       
                     .o    (w36_mabu1     )      
);
DSPCELL_SELBUF #(36) U_DSPCELL_SELBUF_U2(  //assign o = sel == 0 ? o_buf :  i
                     .clk  (clk_mult_u           ),       
                     .rst_n(rst_n         ),       
                     .i    (w36_mabu1     ),     
                     .sel  (cfg_mult_u[1] ),       
                     .o    (w36_mabu2     )    
);
//DSPCELL_MUX2 #(36) U_DSPCELL_MUX2_U3(
//                .i0   (w36_mabu2 ),
//                .i1   (36'h0     ),
//                .sel  (MCTRL[1]  ),
//                .o    (w36_mabu3 )
//);
DSPCELL_MUX2 #(36) U_DSPCELL_MUX2_U3(
                .i0   (36'h0 	 ),
                .i1   (w36_mabu2 ),
                .sel  (MCTRL[1]  ),
                .o    (w36_mabu3 )
);
//DSPCELL_MUX2 #(53) U_DSPCELL_MUX2_U4(
//                .i0   ({w36_mabu3,17'h0}            ),
//                .i1   ({{17{w36_mabu3[35]}},w36_mabu3} ),
//                .sel  (MCTRL[2]                     ),
//                .o    (w53_mabu4                    )
//);
//DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_U5(
//                .i0   ({{3{w53_mabu4[52]}},w53_mabu4}      ),
//                .i1   (U_buf                            ),
//                .sel  (MCTRL[3]                     ),
//                .o    (MR_U                         )
//);
DSPCELL_MUX4 #(56) U_DSPCELL_MUX4_U5(
                .i0   ({{3{w36_mabu3[35]}},w36_mabu3,17'h0}            ),
                .i1   ({{20{w36_mabu3[35]}},w36_mabu3} ),
                .i2   ({{4{w36_mabu3[35]}},w36_mabu3,16'h0}            ),
                .i3   (U_buf                            ),
                .sel  (MCTRL[3:2]                   ),
                .o    (MR_U                         )
);



//=============================================
DSPCELL_MULT #(18) U_DSPCELL_MULT_MABL(
                     .i0 (MA_L      ),
                     .i1 (MB_L      ),
                     .o  (w36_mabl  ) 
);
DSPCELL_SELBUF #(36) U_DSPCELL_SELBUF_L1(  //assign o = sel == 0 ? o_buf :  i
                     .clk  (clk_mult_l           ),       
                     .rst_n(rst_n         ),
                     .i    (w36_mabl      ),     
                     .sel  (cfg_mult_l[0] ),       
                     .o    (w36_mabl1     )      
);
DSPCELL_SELBUF #(36) U_DSPCELL_SELBUF_L2(  //assign o = sel == 0 ? o_buf :  i
                     .clk  (clk_mult_l           ),       
                     .rst_n(rst_n         ),
                     .i    (w36_mabl1     ),     
                     .sel  (cfg_mult_l[1] ),       
                     .o    (w36_mabl2     )    
);
//DSPCELL_MUX2 #(36) U_DSPCELL_MUX2_L3(
//                .i0   (w36_mabl2 ),
//                .i1   (36'h0     ),
//                .sel  (MCTRL[0]  ),
//                .o    (w36_mabl3 )
//);
DSPCELL_MUX2 #(36) U_DSPCELL_MUX2_L3(
                .i0   (36'h0 	 ),
                .i1   (w36_mabl2 ),
                .sel  (MCTRL[0]  ),
                .o    (w36_mabl3 )
);
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_L4(
                .i0   ({{20{w36_mabl3[35]}},w36_mabl3} ),
                .i1   (w56_mcat    ),
                .sel  (MCTRL[4]                     ),
                .o    (MR_L_t                         )
);
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_L5(
                .i0   (MR_L_t),
                .i1   (R[55:0]),
                .sel  (MCTRL[5]                     ),
                .o    (MR_L                         )
);


assign  w56_mcat = {MA_U[1:0],MB_U[17:0],MB_L[17:0],MA_L[17:0]};



endmodule
//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_postadder(
                        clk_poa             ,                  
                        rst_n           ,                    
                        MR_U            ,                   
                        MR_L            ,                   
                        UFC             ,                   
                        R_CARRY_CAS_IN  ,                              
                        R_CARRY_CAS_OUT ,                              
                        R_ECARRY_CAS_IN  ,                              
                        R_ECARRY_CAS_OUT ,                              
                        R_pre           ,                    
                        R               ,                    
                        R_CAS_OUT       ,
                        MATCH           ,
                        RNDM            ,                      
                        SUBCTRL         ,                      
                        ALUCTRL         ,                      
                        FRCTRL          ,                      
                        CCTRL           ,                      
                        cfg_mat_clr     ,
                        cfg_poa_cyout   ,                            
                        cfg_poa_ceyout  ,                            
                        cfg_poa_ceyin   ,                            
                        cfg_poa_rout                                 
                  );

 

//clock and reset
input           clk_poa;
input           rst_n;   //sys reset

input    [55:0]  MR_U;               // 56  I MultBlock MultBlock calculate result
input    [55:0]  MR_L;               // 56  I MultBlock MultBlock calculate result
input    [55:0]  UFC ;               // 56  I UFCMux  UFC Mux select result
input            R_CARRY_CAS_IN ;    // 1   I Input Carry cascade in
output           R_CARRY_CAS_OUT;    // 1   O Output  Carry cascade out
input            R_ECARRY_CAS_IN ;    // 1   I Input Carry cascade in
output           R_ECARRY_CAS_OUT;    // 1   O Output  Carry cascade out
output   [55:0]  R_pre;              // 56  O R output before buffer and mux, to CompUnit
output   [71:0]  R    ;              // 56  O MAC calculate Output
output   [55:0]  R_CAS_OUT    ;      // 
input            MATCH;
input            RNDM   ;            // 1   I Input Round Control
input    [2:0]   SUBCTRL;            // 3   I Postadder Select and Control to perform Subtraction in post stage operation 
input    [2:0]   ALUCTRL;            // 2   I Postadder Control the functionality of ALU operation 
input    [1:0]   FRCTRL ;            // 2   I Postadder Select final result source 
input    [2:0]   CCTRL  ;            // 3   I Postadder Select the source for rounding method, and perform R_CARRY_CAS_IN and user defined CARRY logic 
        
input            cfg_mat_clr     ;
input            cfg_poa_cyout;      // 1   I Input   cfgmem,postadder carry out control
input           cfg_poa_ceyout;    
input            cfg_poa_ceyin;    
input    [1:0]   cfg_poa_rout ;      // 2   I Input   cfgmem,postadder R out control
        
//======================================      
reg         R_S_55_reg;
wire        w1_poa0;
wire        w1_poa1;
wire [56:0] w57_poa2;
wire [55:0] w56_poa3;
wire [71:0] w56_poa4;
reg  [71:0] w56_poa4_reg;
wire [55:0] w56_poa5;
wire        carry;
wire [55:0] A;
wire [55:0] B;
wire [55:0] U;
wire [55:0] S;
wire [55:0] C;
wire [55:0] R_S;
wire [55:0] MR_U_temp; 

always @(posedge clk_poa or negedge rst_n) begin
    if(rst_n == 0) begin
         R_S_55_reg <= `DLY 1'b0;
    end
    else begin
         R_S_55_reg <= `DLY R_S[55];
    end
end
DSPCELL_MUX4 #(1) U_PostAdder_Mux_PO0(
                          .i0  (1'h0         ),     
                          .i1  (R_S_55_reg    ),     
                          .i2  (MR_L[55]      ),     
                          .i3  (MR_U[55]      ),     
                          .sel (CCTRL[2:1]    ),      
                          .o   (w1_poa0       )  
);
//DSPCELL_MUX2 #(1) U_PostAdder_Mux_PO1(
//                          .i0  (R_CARRY_CAS_IN),
//                          .i1  (RNDM          ),     
//                          .sel (CCTRL[0]    ),      
//                          .o   (w1_poa1       )  
//);
DSPCELL_MUX2 #(1) U_PostAdder_Mux_PO1(
                          .i0  (RNDM		),
                          .i1  (R_CARRY_CAS_IN 	),     
                          .sel (CCTRL[0]    ),      
                          .o   (w1_poa1       )  
);
assign carry = w1_poa0 ^ w1_poa1;
//input            R_ECARRY_CAS_IN ;    // 1   I Input Carry cascade in
//output           R_ECARRY_CAS_OUT;    // 1   O Output  Carry cascade out
//wire      [55:0] MR_U_temp; 
DSPCELL_ADD #(57) U_DSPCELL_ADD_PO2(  //s = i0 + i1
                          .i0  ({1'b0,S[55:0]}    ), 
                          .i1  ({C[55:0],carry}   ), 
                          .s   (w57_poa2          ),
                          .c   (R_ECARRY_CAS_OUT_t  ) 
);
DSPCELL_SELBUF U_DSPCELL_SELBUF_PO3E (  //assign o = sel == 0 ? o_buf :  i
                          .clk       (clk_poa            ),
                          .rst_n     (rst_n          ),  
                          .i         (R_ECARRY_CAS_OUT_t   ),
                          .sel       (cfg_poa_ceyout  ),
                          .o         (R_ECARRY_CAS_OUT) 
);
assign R_S = w57_poa2[55:0];
DSPCELL_SELBUF U_DSPCELL_SELBUF_PO3(  //assign o = sel == 0 ? o_buf :  i
                          .clk       (clk_poa            ),
                          .rst_n     (rst_n          ),  
                          .i         (w57_poa2[56]    ),
                          .sel       (cfg_poa_cyout  ),
                          .o         (R_CARRY_CAS_OUT) 
);

//######################
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_PO4E(
                          .i0  (MR_U                         ),
                          .i1  ({54'h0,R_ECARRY_CAS_IN,1'b0} ),     
                          .sel (cfg_poa_ceyin                ),        
                          .o   (MR_U_temp                    )  
);

DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_PO4(
                          .i0  (MR_U_temp   ),
                          .i1  (~MR_U_temp  ),     
                          .sel (SUBCTRL[2]  ),      
                          .o   (A           )  
);
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_PO5(
                          .i0  (MR_L        ),
                          .i1  (~MR_L       ),     
                          .sel (SUBCTRL[1]  ),      
                          .o   (B           )  
);
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_PO6(
                          .i0  (UFC         ),
                          .i1  (~UFC        ),     
                          .sel (SUBCTRL[0]  ),      
                          .o   (U           )  
);
DSPCELL_BIT_ADD #(56) U_DSPCELL_BIT_ADD_PO7 (
                          .i0  (A  ),
                          .i1  (B  ),
                          .i2  (U  ),
                          .s   (S  ),
                          .c   (C  )  
);
DSPCELL_MUX4 #(56) U_DSPCELL_MUX4_PO8(
                          .i0  (R_S         ),
                          .i1  (S           ),     
                          .i2  (C           ),     
                          .i3  (56'h0       ),     
                          .sel (ALUCTRL[1:0]),      
                          .o   (w56_poa3    )  
);
wire [55:0] w56_poa3_mux;
wire        w1_poa3_sel;
assign      w1_poa3_sel = MATCH && cfg_mat_clr;
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_PO9E(
                          .i0  (w56_poa3    ),
                          .i1  (56'h0       ),     
                          .sel (w1_poa3_sel ),      
                          .o   (w56_poa3_mux )  
);

DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_PO9(
                          .i0  (w56_poa3_mux    ),
                          .i1  (~w56_poa3_mux   ),     
                          .sel (ALUCTRL[2]  ),      
                          .o   (R_pre       )  
);
//DSPCELL_SELBUF #(56)  U_DSPCELL_SELBUF_PO10 (  //assign o = sel == 0 ? o_buf :  i
//                     .clk      (clk_poa              ),
//                     .rst_n    (rst_n            ),  
//                     .i        (R_pre            ),
//                     .sel      (cfg_poa_rout[0]  ),
//                     .o        (w56_poa4         ) 
//);
//DSPCELL_SELBUF #(56)  U_DSPCELL_SELBUF_PO11 (  //assign o = sel == 0 ? o_buf :  i
//                     .clk      (clk_poa                    ),
//                     .rst_n    (rst_n                  ),  
//                     .i        ({MR_U[27:0],MR_L[27:0]} ),
//                     .sel      (cfg_poa_rout[1]  ),
//                     .o        (w56_poa5         ) 
//);
//DSPCELL_MUX4 #(56) U_DSPCELL_MUX4_PO12(
//                          .i0  (R_pre         ),
//                          .i1  (MR_L          ),     
//                          .i2  ({MR_U[27:0],MR_L[27:0]}  ),     
//                          .i3  (56'h0         ),     
//                          .sel (FRCTRL[1:0]   ), 
//                          .o   (w56_poa4      )  
//);
DSPCELL_MUX2 #(72) U_DSPCELL_MUX2_PO10(
                          .i0  ({{16{R_pre[55]}},R_pre}  ),
                          .i1  ({MR_U[35:0],MR_L[35:0]}),     
                          .sel (FRCTRL[0]   ), 
                          .o   (w56_poa4      )  
);
//DSPCELL_SELBUF #(56)  U_DSPCELL_SELBUF_PO10 (  //assign o = sel == 0 ? o_buf :  i
//                     .clk      (clk_poa              ),
//                     .rst_n    (rst_n            ),  
//                     .i        (w56_poa4 ),
//                     .sel      (cfg_poa_rout[0]  ),
//                     .o        (R         ) 
//);
always @(posedge clk_poa or negedge rst_n) begin
    if(rst_n == 0) begin
         w56_poa4_reg <= 56'b0;
    end
    else begin
         w56_poa4_reg <= w56_poa4;
    end
end
DSPCELL_MUX2 #(72)  U_DSPCELL_MUX2_PO11 (
                     .i0       	(w56_poa4_reg 	),
		     .i1	(w56_poa4	),
                     .sel      	(cfg_poa_rout[0]),
                     .o        	(R         ) 
);
//DSPCELL_SELBUF #(56)  U_DSPCELL_SELBUF_PO11 (  //assign o = sel == 0 ? o_buf :  i
//                     .clk      (clk_poa                    ),
//                     .rst_n    (rst_n                  ),  
//                     .i        (w56_poa4 ),
//                     .sel      (cfg_poa_rout[1]  ),
//                     .o        (R_CAS_OUT         ) 
//);
DSPCELL_MUX2 #(56)  U_DSPCELL_MUX2_PO12 (
                     .i0        (w56_poa4_reg[55:0] ),
		     .i1	(w56_poa4[55:0]	    ),
                     .sel      	(cfg_poa_rout[1]    ),
                     .o        	(R_CAS_OUT         ) 
);


endmodule
//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_preadder(
                      clk_pra          ,                     
                      rst_n        ,
                      A_L          ,                     
                      C_L          ,                     
                      D_L          ,                     
                      A_U          ,                     
                      C_U          ,                     
                      D_U          ,                     
                      A_L_CAS_IN   ,                            
                      C_L_CAS_IN   ,                            
                      A_U_CAS_IN   ,                            
                      C_U_CAS_IN   ,                            
                      A_L_CAS_OUT  ,                             
                      C_L_CAS_OUT  ,                             
                      A_U_CAS_OUT  ,                             
                      C_U_CAS_OUT  ,                             
                      MA_U         ,   
                      MB_U         ,   
                      MB_L         ,   
                      MA_L         ,   
                      PAZCTRL      ,    
                      PARCTRL      ,    
                      PASUBCTRL    ,      
                      BLCTRL       ,                        
                      BUCTRL       ,                        
                      PASCTRL      ,    
                      cfg_pra_au   ,                            
                      cfg_pra_cu   ,                            
                      cfg_pra_du   ,                            
                      cfg_pra_dl   ,                            
                      cfg_pra_al   ,                            
                      cfg_pra_cl   ,                            
                      cfg_pra_ou   ,                                                           
                      cfg_pra_ol                                
                  );

 

//clock and reset
input           clk_pra;
input           rst_n;   //sys reset

input  [17:0]   A_L;            //Input Input of the lower multiplier 
input  [17:0]   C_L;            //Input Input to the Pre-Adder and can be used as another input to the lower multiplier 
input  [17:0]   D_L;            //Input Another input to the Pre-Adder 
input  [17:0]   A_U;            //Input Input of the upper multiplier 
input  [17:0]   C_U;            //Input Input to the Pre-Adder and can be used as another input to the upper multiplier 
input  [17:0]   D_U;            //Input Another input to the Pre-Adder 
        
input  [17:0]   A_L_CAS_IN;     //Input Cascaded data input from A_L_CAS_OUT of previous DSP slice 
input  [17:0]   C_L_CAS_IN;     //Input Cascaded data input from C_L_CAS_OUT of previous DSP slice 
input  [17:0]   A_U_CAS_IN;     //Input Cascaded data input from A_U_CAS_OUT of previous DSP slice 
input  [17:0]   C_U_CAS_IN;     //Input Cascaded data input from C_U_CAS_OUT of previous DSP slice 
        
output [17:0]   A_L_CAS_OUT;    //Output  Cascaded data output to A_L_CAS_IN of next DSP slice 
output [17:0]   C_L_CAS_OUT;    //Output  Cascaded data output to C_L_CAS_IN of next DSP slice 
output [17:0]   A_U_CAS_OUT;    //Output  Cascaded data output to A_U_CAS_IN of next DSP slice 
output [17:0]   C_U_CAS_OUT;    //Output  Cascaded data output to C_U_CAS_IN of next DSP slice 

output [17:0]   MA_U;   
output [17:0]   MB_U;   
output [17:0]   MB_L;   
output [17:0]   MA_L;   
        
                                //Select and Control the functionality of the Pre-Adder and Selector
input  [5:0]    PAZCTRL; 
input  [5:0]    PARCTRL; 
input  [1:0]    PASUBCTRL; 
input           BLCTRL; 
input           BUCTRL; 
input  [7:0]    PASCTRL;

input  [2:0]    cfg_pra_au;     //3 I Input cfg mempreadder AU control
input  [2:0]    cfg_pra_cu;     //3 I Input cfg mempreadder CU control
input           cfg_pra_du;     //1 I Input cfg mempreadder DU control
input           cfg_pra_dl;     //1 I Input cfg mempreadder DL control
input  [2:0]    cfg_pra_al;     //3 I Input cfg mempreadder AL control
input  [2:0]    cfg_pra_cl;     //3 I Input cfg mempreadder CL control
input           cfg_pra_ou;     //1 I Input cfg mempreadder OU control
input           cfg_pra_ol;     //1 I Input cfg mempreadder OL control

wire   [17:0]   w18_au0;
wire   [17:0]   w18_au1;
wire   [17:0]   w18_au2;
wire   [17:0]   w18_au3;
wire   [17:0]   w18_cu0;
wire   [17:0]   w18_cu1;
wire   [17:0]   w18_cu2;
wire   [17:0]   w18_cu3;
wire   [17:0]   w18_du2;
wire   [17:0]   w18_du3;
wire   [17:0]   w18_dl2;
wire   [17:0]   w18_dl3;
wire   [17:0]   w18_cl0;
wire   [17:0]   w18_cl1;
wire   [17:0]   w18_cl2;
wire   [17:0]   w18_cl3;
wire   [17:0]   w18_al0;
wire   [17:0]   w18_al1;
wire   [17:0]   w18_al2;
wire   [17:0]   w18_al3;

wire   [17:0]   D_U_CAS_OUT;    //Output  Cascaded data output to A_U_CAS_IN of next DSP slice 
wire   [17:0]   D_L_CAS_OUT;    //Output  Cascaded data output to C_U_CAS_IN of next DSP slice 
wire   [17:0]   A_U_BP;
wire   [17:0]   B_U;
wire   [17:0]   A_L_BP;
wire   [17:0]   B_L;
wire   [17:0]   w18_bu_0;
wire   [17:0]   w18_bu_1;
wire   [17:0]   w18_bu_2;
wire   [17:0]   w18_bu_3;
wire   [17:0]   w18_bl_0;
wire   [17:0]   w18_bl_1;
wire   [17:0]   w18_bl_2;
wire   [17:0]   w18_bl_3;
wire   [17:0]   C_U_CAS_OUT_t;
wire   [17:0]   C_L_CAS_OUT_t;

//======================================      
//AU 5
DSPCELL_MUX2 #(18) U_PAMUX_AU0(
                          .i0  (A_L_CAS_OUT   ),     
                          .i1  (A_U_CAS_IN    ),     
                          .sel (cfg_pra_au[0] ),      
                          .o   (w18_au0         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_AU1(
                          .i0  (w18_au0         ),     
                          .i1  (A_U           ),     
                          .sel (cfg_pra_au[1] ),      
                          .o   (w18_au1         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_AU2(
                          .i0  (18'h0           ),     
                          .i1  (w18_au1         ),     
                          .sel (PAZCTRL[5]      ),      
                          .o   (w18_au2         )  
);

//DSPCELL_AND2 #(18) U_PAAND2_AU2(
//                          .i0  (PAZCTRL[5]    ),
//                          .i1  (w18_au1         ),
//                          .o   (w18_au2         )
//);

DSPCELL_SELBUF #(18) U_PCELL_SELBUF_AU3(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_au2         ),  
                          .sel (cfg_pra_au[2] ),   
                          .o   (w18_au3         ) 
);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_AU4(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_au3         ),  
                          .sel (PARCTRL[5]    ),   
                          .o   (A_U_CAS_OUT   ) 
);

//CU 4
DSPCELL_MUX2 #(18) U_PAMUX_CU0(
                          .i0  (C_L_CAS_OUT   ),     
                          .i1  (C_U_CAS_IN    ),     
                          .sel (cfg_pra_cu[0] ),      
                          .o   (w18_cu0         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_CU1(
                          .i0  (w18_cu0         ),     
                          .i1  (C_U           ),     
                          .sel (cfg_pra_cu[1] ),      
                          .o   (w18_cu1         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_CU2(
                          .i0  (18'h0           ),     
                          .i1  (w18_cu1         ),     
                          .sel (PAZCTRL[4]      ),      
                          .o   (w18_cu2         )  
);

//
//DSPCELL_AND2 #(18) U_PAAND2_CU2(
//                          .i0  (PAZCTRL[4]    ),
//                          .i1  (w18_cu1         ),
//                          .o   (w18_cu2         )
//);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_CU3(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_cu2         ),  
                          .sel (cfg_pra_cu[2] ),   
                          .o   (w18_cu3         ) 
);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_CU4(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_cu3         ),  
                          .sel (PARCTRL[4]    ),   
                          .o   (C_U_CAS_OUT   ) 
);
DSPCELL_MUX2 #(18)  U_PAMUX_BU0(
                          .i0  (C_U_CAS_OUT   ), 
                          .i1  (~C_U_CAS_OUT  ),
                          .sel (PASUBCTRL[1]  ),      
                          .o   (C_U_CAS_OUT_t )  
);

//DU 3
DSPCELL_MUX2 #(18) U_PAMUX_DU2(
                          .i0  (18'h0           ),     
                          .i1  (D_U             ),     
                          .sel (PAZCTRL[3]      ),      
                          .o   (w18_du2         )  
);
//DSPCELL_AND2 #(18) U_PAAND2_DU2(
//                          .i0  (PAZCTRL[3]    ),
//                          .i1  (D_U           ),
//                          .o   (w18_du2         )
//);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_DU3(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_du2         ),  
                          .sel (cfg_pra_du    ),   
                          .o   (w18_du3         ) 
);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_DU4(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_du3         ),  
                          .sel (PARCTRL[3]    ),   
                          .o   (D_U_CAS_OUT   ) 
);

//DL 2
DSPCELL_MUX2 #(18) U_PAMUX_DL2(
                          .i0  (18'h0           ),     
                          .i1  (D_L             ),     
                          .sel (PAZCTRL[2]      ),      
                          .o   (w18_dl2         )  
);

//DSPCELL_AND2 #(18) U_PAAND2_DL2(
//                          .i0  (PAZCTRL[2]    ),
//                          .i1  (D_L           ),
//                          .o   (w18_dl2         )
//);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_DL3(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_dl2         ),  
                          .sel (cfg_pra_dl    ),   
                          .o   (w18_dl3         ) 
);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_DL4(
                          .clk (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i   (w18_dl3         ),  
                          .sel (PARCTRL[2]    ),   
                          .o   (D_L_CAS_OUT   ) 
);


//CL 1
DSPCELL_MUX2 #(18) U_PAMUX_CL0(
                          .i0  (C_L_CAS_IN    ),     
                          .i1  (C_U_CAS_IN    ),     
                          .sel (cfg_pra_cl[0] ),      
                          .o   (w18_cl0         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_CL1(
                          .i0  (w18_cl0         ),     
                          .i1  (C_L           ),     
                          .sel (cfg_pra_cl[1] ),      
                          .o   (w18_cl1         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_CL2(
                          .i0  (18'h0           ),     
                          .i1  (w18_cl1         ),     
                          .sel (PAZCTRL[1]      ),      
                          .o   (w18_cl2         )  
);


//DSPCELL_AND2 #(18) U_PAAND2_CL2(
//                          .i0  (PAZCTRL[1]    ),
//                          .i1  (w18_cl1         ),
//                          .o   (w18_cl2         )
//);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_CL3(
                          .clk  (clk_pra            ),  
                          .rst_n(rst_n          ),       
                          .i    (w18_cl2        ),  
                          .sel  (cfg_pra_cl[2]  ),   
                          .o    (w18_cl3        ) 
);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_CL4(
                          .clk  (clk_pra            ),  
                          .rst_n(rst_n          ),       
                          .i    (w18_cl3        ),  
                          .sel  (PARCTRL[1]     ),   
                          .o    (C_L_CAS_OUT    ) 
);
DSPCELL_MUX2 #(18)  U_PAMUX_BL0(
                          .i0  (C_L_CAS_OUT   ), 
                          .i1  (~C_L_CAS_OUT  ),
                          .sel (PASUBCTRL[0]  ),      
                          .o   (C_L_CAS_OUT_t )  
);
//AL 0
DSPCELL_MUX2 #(18) U_PAMUX_AL0(
                          .i0  (A_L_CAS_IN      ),     
                          .i1  (A_U_CAS_IN      ),     
                          .sel (cfg_pra_al[0]   ),      
                          .o   (w18_al0         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_AL1(
                          .i0  (w18_al0         ),     
                          .i1  (A_L             ),     
                          .sel (cfg_pra_al[1]   ),      
                          .o   (w18_al1         )  
);
DSPCELL_MUX2 #(18) U_PAMUX_AL2(
                          .i0  (18'h0           ),     
                          .i1  (w18_al1         ),     
                          .sel (PAZCTRL[0]      ),      
                          .o   (w18_al2         )  
);

//DSPCELL_AND2 #(18) U_PAAND2_AL2(
//                          .i0  (PAZCTRL[1]      ),
//                          .i1  (w18_al1         ),
//                          .o   (w18_al2         )
//);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_AL3(
                          .clk    (clk_pra           ),  
                          .rst_n  (rst_n         ),       
                          .i      (w18_al2       ),  
                          .sel    (cfg_pra_al[2] ),   
                          .o      (w18_al3       ) 
);
DSPCELL_SELBUF #(18) U_PCELL_SELBUF_AL4(
                          .clk    (clk_pra           ),  
                          .rst_n  (rst_n         ),       
                          .i      (w18_al3       ),  
                          .sel    (PARCTRL[0]    ),   
                          .o      (A_L_CAS_OUT   ) 
);

assign A_U_BP = A_U_CAS_OUT;
assign A_L_BP = A_L_CAS_OUT;
//BU
//DSPCELL_MUX2 #(18)  U_PAMUX_BU0(
//                          .i0  (D_U_CAS_OUT   ), 
//                          .i1  (~D_U_CAS_OUT  ),
//                          .sel (PASUBCTRL[1]  ),      
//                          .o   (w18_bu_0      )  
//);
assign w18_bu_0 = D_U_CAS_OUT ;
DSPCELL_FULLADD #(18)   U_PCELL_FULLADD_BU1  (  //s = i0 + i1
                     .i0   (C_U_CAS_OUT_t),
                     .i1   (w18_bu_0     ),
                     .s    (w18_bu_1     ),
                     .ci   (PASUBCTRL[1] ),
                     .co   (             )  
);
DSPCELL_SELBUF #(18)  U_PCELL_SELBUF_BU2(
                          .clk  (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i    (w18_bu_1      ),  
                          .sel  (cfg_pra_ou    ),   
                          .o    (w18_bu_2      ) 
);
DSPCELL_MUX2 #(18)  U_PAMUX_BU3(
                          .i0  (C_U_CAS_OUT ),     
                          .i1  (w18_bu_2      ),     
                          .sel (BUCTRL        ),      
                          .o   (B_U           )  
);
//BL
//DSPCELL_MUX2 #(18)  U_PAMUX_BL0(
//                          .i0  (D_L_CAS_OUT   ), 
//                          .i1  (~D_L_CAS_OUT  ),
//                          .sel (PASUBCTRL[0]  ),      
//                          .o   (w18_bl_0      )  
//);
assign w18_bl_0 = D_L_CAS_OUT ;
DSPCELL_FULLADD #(18)   U_PCELL_FULLADD_BL1  (  //s = i0 + i1
                     .i0   (C_L_CAS_OUT_t),
                     .i1   (w18_bl_0     ),
                     .s    (w18_bl_1     ),
                     .ci   (PASUBCTRL[0] ),
                     .co   (             )  
);
DSPCELL_SELBUF #(18)  U_PCELL_SELBUF_BL2(
                          .clk  (clk_pra           ),  
                          .rst_n(rst_n         ),       
                          .i    (w18_bl_1      ),  
                          .sel  (cfg_pra_ol    ),   
                          .o    (w18_bl_2      ) 
);
DSPCELL_MUX2 #(18)  U_PAMUX_BL4(
                          .i0  (C_L_CAS_OUT ),     
                          .i1  (w18_bl_2      ),     
                          .sel (BLCTRL        ),      
                          .o   (B_L           )  
);
//BL
//PCELL_ADD #(18)   U_PCELL_ADD_BL0  (  //s = i0 + i1
//                     .i0   (C_L_CAS_OUT  ),
//                     .i1   (D_L_CAS_OUT  ),
//                     .s    (w18_bl_0     ),
//                     .c    (             )  
//);
//DSPCELL_SUB #(18) U_DSPCELL_SUB_BL1  (  // s = i0 - i1
//                     .i0   (C_L_CAS_OUT  ),
//                     .i1   (D_L_CAS_OUT  ),
//                     .s    (w18_bl_1     ),
//                     .c    (             ) 
//);
//DSPCELL_MUX2 #(18)  U_PAMUX_BL2(
//                          .i0  (w18_bl_0      ), //add 
//                          .i1  (w18_bl_1      ), //sub  
//                          .sel (PASUBCTRL[0]  ),      
//                          .o   (w18_bl_2      )  
//);
//PCELL_SELBUF #(18)  U_PCELL_SELBUF_BL3(
//                          .clk  (clk           ),  
//                          .rst_n(rst_n         ),       
//                          .i    (w18_bl_2      ),  
//                          .sel  (cfg_pra_ol    ),   
//                          .o    (w18_bl_3      ) 
//);
//DSPCELL_MUX2 #(18)  U_PAMUX_BL4(
//                          .i0  (C_U_CAS_OUT   ),     
//                          .i1  (w18_bl_3      ),     
//                          .sel (BLCTRL        ),
//                          .o   (B_L           )  
//);
//MA_U
DSPCELL_MUX4 #(18) U_DSPCELL_MUX4_MA_U(
                     .i3   (A_U_BP       ),  
                     .i2   (B_U          ),  
                     .i1   (A_L_BP       ),  
                     .i0   (B_L          ),  
                     .sel  (PASCTRL[7:6] ),   
                     .o    (MA_U         ) 
);
//MB_U
DSPCELL_MUX4 #(18) U_DSPCELL_MUX4_MB_U(
                     .i3   (A_U_BP       ),  
                     .i2   (B_U          ),  
                     .i1   (A_L_BP       ),  
                     .i0   (B_L          ),  
                     .sel  (PASCTRL[5:4] ),   
                     .o    (MB_U         ) 
);
//MB_L
DSPCELL_MUX4 #(18) U_DSPCELL_MUX4_MB_L(
                     .i3   (A_U_BP       ),  
                     .i2   (B_U          ),  
                     .i1   (A_L_BP       ),  
                     .i0   (B_L          ),  
                     .sel  (PASCTRL[3:2] ),   
                     .o    (MB_L         ) 
);
//MA_L
DSPCELL_MUX4 #(18) U_DSPCELL_MUX4_MA_L(
                     .i3   (A_U_BP       ),  
                     .i2   (B_U          ),  
                     .i1   (A_L_BP       ),  
                     .i0   (B_L          ),  
                     .sel  (PASCTRL[1:0] ),   
                     .o    (MA_L         ) 
);

endmodule
//*************************************************
//company:   capital-micro
//author:   hongyu.wang
//date:      20140526
//function:   `DSP
//*************************************************
//$Log: .v,v $


`ifndef DLY
`define DLY #0.1
`endif


module dsp_ufcmux(
                   clk_ufc          ,    
                   rst_n        ,
                   R_CAS_IN     ,           
                   R            ,    
                   U            ,    
                   UFC          ,      
                   U_BUF        ,        
                   FCCTRL       ,       
                   UFCCTRL      ,        
                   cfg_ufcmux               
                                     );
//clock and reset
input           clk_ufc;
input           rst_n;   //sys reset

input  [55:0]   R_CAS_IN;  
input  [55:0]   R;  
input  [55:0]   U;  
output [55:0]   UFC;  
output [55:0]   U_BUF;  

input  [2:0]    FCCTRL;
input           UFCCTRL;
input           cfg_ufcmux;

reg    [55:0]   R_CAS_IN_buf;
wire   [55:0]   w56_ufcmux0;

always @(posedge clk_ufc or negedge rst_n ) begin
    if(rst_n == 0) begin
        R_CAS_IN_buf <= `DLY 56'h0;
    end
    else begin
        R_CAS_IN_buf <= `DLY R_CAS_IN;
    end
end
//DSPCELL_MUX8 #(56) U_PCELL_MUX8_UFCMUX0(
//                     .i0  ( R                                   ), 
//                     .i1  ( 56'h0                               ), 
//                     .i2  ( {{17{R[55]}},R[55:17]}                ), 
//                     .i3  ( {{34{R[55]}},R[55:34]}                ), 
//                     .i4  ( R_CAS_IN                            ), 
//                     .i5  ( {{34{R_CAS_IN[55]}},R_CAS_IN[55:34]}  ), 
//                     .i6  ( R_CAS_IN_buf                        ), 
//                     .i7  ( {{17{R_CAS_IN[55]}},R_CAS_IN[55:17]}  ), 
//                     .sel ( FCCTRL                              ),  
//                     .o   ( w56_ufcmux0                         )  
//);
DSPCELL_MUX8 #(56) U_PCELL_MUX8_UFCMUX0(
                     .i0  ( 56'h0                                   ), 
                     .i1  ( R                               ), 
                     .i2  ( {{17{R[55]}},R[55:17]}                ), 
                     .i3  ( {{34{R[55]}},R[55:34]}                ), 
                     .i4  ( R_CAS_IN                            ), 
                     .i5  ( {{34{R_CAS_IN[55]}},R_CAS_IN[55:34]}  ), 
                     .i6  ( R_CAS_IN_buf                        ), 
                     .i7  ( {{17{R_CAS_IN[55]}},R_CAS_IN[55:17]}  ), 
                     .sel ( FCCTRL                              ),  
                     .o   ( w56_ufcmux0                         )  
);

DSPCELL_SELBUF #(56) U_PCELL_SELBUF_UFCMUX1(  //assign o = sel == 0 ? o_buf :  i
                     .clk ( clk_ufc         ),    
                     .rst_n ( rst_n),    
                     .i   ( U           ),  
                     .sel ( cfg_ufcmux  ),    
                     .o   ( U_BUF       )   
);
//DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_UFCMUX2(
//                .i0   (U_BUF           ),
//                .i1   (w56_ufcmux0     ),
//                .sel  (UFCCTRL         ),
//                .o    (UFC             )
//);
DSPCELL_MUX2 #(56) U_DSPCELL_MUX2_UFCMUX2(
                .i0   (w56_ufcmux0     ),
                .i1   (U_BUF           ),
                .sel  (UFCCTRL         ),
                .o    (UFC             )
);

endmodule
//================================================================================
// Copyright (c) 2012 Capital-micro, Inc.(Beijing)  All rights reserved.
//
// Capital-micro, Inc.(Beijing) Confidential.
//
// No part of this code may be reproduced, distributed, transmitted,
// transcribed, stored in a retrieval system, or translated into any
// human or computer language, in any form or by any means, electronic,
// mechanical, magnetic, manual, or otherwise, without the express
// written permission of Capital-micro, Inc.
//
//================================================================================
// Module Description: 
// This is the decoder module of the ECC IP 
//================================================================================
// Revision History :
//     V1.0   2012-11-30  FPGA IP Grp, first created
//     V1.1   2012-12-03  FPGA IP Grp, Add pipeline_en for timing performance
//================================================================================
module ECC_DECODER(
    i_data,
    i_parity,
    eccoutdberr,
    eccoutsberr,
    o_code,
    o_parity
);

//---------------------------------------------------------------------
// inputs & outputs
//---------------------------------------------------------------------
input   [63:0]  i_data;
input   [7:0]   i_parity;
output  eccoutdberr;
output  eccoutsberr;
output  [63:0]  o_code;
output  [7:0] o_parity;

wire [71:0] data_wire;
wire [63:0] code_wire;
wire [7:0] parity_wire;

assign data_wire = {i_data[63:57],i_parity[7],i_data[56:26],i_parity[6],i_data[25:11],i_parity[5],i_data[10:4],i_parity[4],i_data[3:1],i_parity[3],
                      i_data[0],i_parity[2:0]};

assign o_parity	    = parity_wire;
assign o_code	    = code_wire;

//---------------------------------------------------------------------
// instantiate module
//---------------------------------------------------------------------
ecc_decoder_core inst_ecc_decoder_core(
    .i_data             (data_wire),
    .o_err_corrected    (eccoutsberr),
    .o_err_fatal        (eccoutdberr),
    .o_code             (code_wire),
    .o_parity		(parity_wire)
);

endmodule


//---------------------------------------------------------------------
// Core ECC decoder module
//---------------------------------------------------------------------
module ecc_decoder_core(
    i_data,
    o_err_corrected,
    o_err_fatal,
    o_code,
    o_parity
);
localparam data_width = 72;
localparam parity_width = (data_width > 15 && data_width <= 31 ) ? 6 :
                          (data_width > 31 && data_width <= 63 ) ? 7 :
                          (data_width > 63 && data_width <= 127) ? 8 :
                          0; // 0 means not support

localparam code_width = data_width - parity_width;
localparam error_bit_width = 1 << (parity_width - 1);

input   [(data_width)-1:0]  i_data;
output                      o_err_corrected;
output                      o_err_fatal;
output  [(code_width)-1:0]  o_code;
output  [(parity_width)-1:0] o_parity;

wire [(parity_width)-1:0]   syndrome;
wire [(data_width)-1:0]     x;
wire syndrome_err;
wire parity_err;
wire data_err;
wire [(error_bit_width)-1:0]error_bit;
wire [(code_width)-1:0]     x_data_wire;
wire [(parity_width)-1:0]   x_parity_wire;
wire [(parity_width)-1:0]   syndrome_wire;

reg [(code_width)-1:0]      x_data_r;
reg [(parity_width)-1:0]    x_parity_r;
reg [(parity_width)-1:0]    syndrome_r;

assign x = i_data;
assign o_err_corrected = syndrome_wire[0];                                  //only-1-error-occuring and corrected
assign o_err_fatal     = syndrome_err & (~(syndrome_wire[0])) ;             //2-errors detected

error_bit_decoder inst_error_bit_decoder(
    .i_data     (syndrome_wire[(parity_width)-1:1]),
    .o_decodes  (error_bit)
);
defparam inst_error_bit_decoder.data_width = parity_width - 1;

        //parity check
        assign syndrome[7]    = x[64]^(^x[71:65]);
        assign syndrome[6]    = x[32]^(^x[63:33]);
        assign syndrome[5]    = x[16]^(^x[63:48])^(^x[31:17]);
        assign syndrome[4]    = x[ 8]^(^x[63:56])^(^x[47:40])^(^x[31:24])^(^x[15:9]);
        assign syndrome[3]    = x[ 4]^(^x[71:68])^(^x[63:60])^(^x[55:52])^(^x[47:44])^(^x[39:36])^(^x[31:28])^(^x[23:20])^(^x[15:12])^(^x[7:5]);
        assign syndrome[2]    = x[ 2]^(^x[71:70])^(^x[67:66])^(^x[63:62])^(^x[59:58])^(^x[55:54])^(^x[51:50])^(^x[47:46])^(^x[43:42])^(^x[39:38])^(^x[35:34])^(^x[31:30])^(^x[27:26])^(^x[23:22])^(^x[19:18])^(^x[15:14])^(^x[11:10])^(^x[7:6])^x[3];
        assign syndrome[1]    = x[ 1]^x[71]^x[69]^x[67]^x[65]^x[63]^x[61]^x[59]^x[57]^x[55]^x[53]^x[51]^x[49]^x[47]^x[45]^x[43]^x[41]^x[39]^x[37]^x[35]^x[33]^x[31]^x[29]^x[27]^x[25]^x[23]^x[21]^x[19]^x[17]^x[15]^x[13]^x[11]^x[9]^x[7]^x[5]^x[3];
        //extra-parity-bit
        assign syndrome[0]    = x[ 0]^(^x[71:1]);

        assign x_data_wire  = {x[71:65],x[63:33],x[31:17],x[15:9],x[7:5],x[3]};
	assign x_parity_wire = {x[64],x[32],x[16],x[8],x[4],x[2],x[1],x[0]}; 
	assign syndrome_wire= syndrome;

        //nonzero/error check
        assign syndrome_err = |syndrome_wire[7:1];
        assign parity_err   = error_bit[64]|error_bit[32]|error_bit[16]|error_bit[8]|error_bit[4]|error_bit[2]|error_bit[1];
        assign data_err     = (|error_bit[71:65])|(|error_bit[63:33])|(|error_bit[31:17])|(|error_bit[15:9])|(|error_bit[7:5])|error_bit[3];
        //output code (corrected when only-1-error-occuring)
        assign o_code[63]   = syndrome_wire[0] ? error_bit[71]^x_data_wire[63] : x_data_wire[63];
        assign o_code[62]   = syndrome_wire[0] ? error_bit[70]^x_data_wire[62] : x_data_wire[62];
        assign o_code[61]   = syndrome_wire[0] ? error_bit[69]^x_data_wire[61] : x_data_wire[61];
        assign o_code[60]   = syndrome_wire[0] ? error_bit[68]^x_data_wire[60] : x_data_wire[60];
        assign o_code[59]   = syndrome_wire[0] ? error_bit[67]^x_data_wire[59] : x_data_wire[59];
        assign o_code[58]   = syndrome_wire[0] ? error_bit[66]^x_data_wire[58] : x_data_wire[58];
        assign o_code[57]   = syndrome_wire[0] ? error_bit[65]^x_data_wire[57] : x_data_wire[57];
        assign o_code[56]   = syndrome_wire[0] ? error_bit[63]^x_data_wire[56] : x_data_wire[56];
        assign o_code[55]   = syndrome_wire[0] ? error_bit[62]^x_data_wire[55] : x_data_wire[55];
        assign o_code[54]   = syndrome_wire[0] ? error_bit[61]^x_data_wire[54] : x_data_wire[54];
        assign o_code[53]   = syndrome_wire[0] ? error_bit[60]^x_data_wire[53] : x_data_wire[53];
        assign o_code[52]   = syndrome_wire[0] ? error_bit[59]^x_data_wire[52] : x_data_wire[52];
        assign o_code[51]   = syndrome_wire[0] ? error_bit[58]^x_data_wire[51] : x_data_wire[51];
        assign o_code[50]   = syndrome_wire[0] ? error_bit[57]^x_data_wire[50] : x_data_wire[50];
        assign o_code[49]   = syndrome_wire[0] ? error_bit[56]^x_data_wire[49] : x_data_wire[49];
        assign o_code[48]   = syndrome_wire[0] ? error_bit[55]^x_data_wire[48] : x_data_wire[48];
        assign o_code[47]   = syndrome_wire[0] ? error_bit[54]^x_data_wire[47] : x_data_wire[47];
        assign o_code[46]   = syndrome_wire[0] ? error_bit[53]^x_data_wire[46] : x_data_wire[46];
        assign o_code[45]   = syndrome_wire[0] ? error_bit[52]^x_data_wire[45] : x_data_wire[45];
        assign o_code[44]   = syndrome_wire[0] ? error_bit[51]^x_data_wire[44] : x_data_wire[44];
        assign o_code[43]   = syndrome_wire[0] ? error_bit[50]^x_data_wire[43] : x_data_wire[43];
        assign o_code[42]   = syndrome_wire[0] ? error_bit[49]^x_data_wire[42] : x_data_wire[42];
        assign o_code[41]   = syndrome_wire[0] ? error_bit[48]^x_data_wire[41] : x_data_wire[41];
        assign o_code[40]   = syndrome_wire[0] ? error_bit[47]^x_data_wire[40] : x_data_wire[40];
        assign o_code[39]   = syndrome_wire[0] ? error_bit[46]^x_data_wire[39] : x_data_wire[39];
        assign o_code[38]   = syndrome_wire[0] ? error_bit[45]^x_data_wire[38] : x_data_wire[38];
        assign o_code[37]   = syndrome_wire[0] ? error_bit[44]^x_data_wire[37] : x_data_wire[37];
        assign o_code[36]   = syndrome_wire[0] ? error_bit[43]^x_data_wire[36] : x_data_wire[36];
        assign o_code[35]   = syndrome_wire[0] ? error_bit[42]^x_data_wire[35] : x_data_wire[35];
        assign o_code[34]   = syndrome_wire[0] ? error_bit[41]^x_data_wire[34] : x_data_wire[34];
        assign o_code[33]   = syndrome_wire[0] ? error_bit[40]^x_data_wire[33] : x_data_wire[33];
        assign o_code[32]   = syndrome_wire[0] ? error_bit[39]^x_data_wire[32] : x_data_wire[32];
        assign o_code[31]   = syndrome_wire[0] ? error_bit[38]^x_data_wire[31] : x_data_wire[31];
        assign o_code[30]   = syndrome_wire[0] ? error_bit[37]^x_data_wire[30] : x_data_wire[30];
        assign o_code[29]   = syndrome_wire[0] ? error_bit[36]^x_data_wire[29] : x_data_wire[29];
        assign o_code[28]   = syndrome_wire[0] ? error_bit[35]^x_data_wire[28] : x_data_wire[28];
        assign o_code[27]   = syndrome_wire[0] ? error_bit[34]^x_data_wire[27] : x_data_wire[27];
        assign o_code[26]   = syndrome_wire[0] ? error_bit[33]^x_data_wire[26] : x_data_wire[26];
        assign o_code[25]   = syndrome_wire[0] ? error_bit[31]^x_data_wire[25] : x_data_wire[25];
        assign o_code[24]   = syndrome_wire[0] ? error_bit[30]^x_data_wire[24] : x_data_wire[24];
        assign o_code[23]   = syndrome_wire[0] ? error_bit[29]^x_data_wire[23] : x_data_wire[23];
        assign o_code[22]   = syndrome_wire[0] ? error_bit[28]^x_data_wire[22] : x_data_wire[22];
        assign o_code[21]   = syndrome_wire[0] ? error_bit[27]^x_data_wire[21] : x_data_wire[21];
        assign o_code[20]   = syndrome_wire[0] ? error_bit[26]^x_data_wire[20] : x_data_wire[20];
        assign o_code[19]   = syndrome_wire[0] ? error_bit[25]^x_data_wire[19] : x_data_wire[19];
        assign o_code[18]   = syndrome_wire[0] ? error_bit[24]^x_data_wire[18] : x_data_wire[18];
        assign o_code[17]   = syndrome_wire[0] ? error_bit[23]^x_data_wire[17] : x_data_wire[17];
        assign o_code[16]   = syndrome_wire[0] ? error_bit[22]^x_data_wire[16] : x_data_wire[16];
        assign o_code[15]   = syndrome_wire[0] ? error_bit[21]^x_data_wire[15] : x_data_wire[15];
        assign o_code[14]   = syndrome_wire[0] ? error_bit[20]^x_data_wire[14] : x_data_wire[14];
        assign o_code[13]   = syndrome_wire[0] ? error_bit[19]^x_data_wire[13] : x_data_wire[13];
        assign o_code[12]   = syndrome_wire[0] ? error_bit[18]^x_data_wire[12] : x_data_wire[12];
        assign o_code[11]   = syndrome_wire[0] ? error_bit[17]^x_data_wire[11] : x_data_wire[11];
        assign o_code[10]   = syndrome_wire[0] ? error_bit[15]^x_data_wire[10] : x_data_wire[10];
        assign o_code[ 9]   = syndrome_wire[0] ? error_bit[14]^x_data_wire[ 9] : x_data_wire[ 9];
        assign o_code[ 8]   = syndrome_wire[0] ? error_bit[13]^x_data_wire[ 8] : x_data_wire[ 8];
        assign o_code[ 7]   = syndrome_wire[0] ? error_bit[12]^x_data_wire[ 7] : x_data_wire[ 7];
        assign o_code[ 6]   = syndrome_wire[0] ? error_bit[11]^x_data_wire[ 6] : x_data_wire[ 6];
        assign o_code[ 5]   = syndrome_wire[0] ? error_bit[10]^x_data_wire[ 5] : x_data_wire[ 5];
        assign o_code[ 4]   = syndrome_wire[0] ? error_bit[ 9]^x_data_wire[ 4] : x_data_wire[ 4];
        assign o_code[ 3]   = syndrome_wire[0] ? error_bit[ 7]^x_data_wire[ 3] : x_data_wire[ 3];
        assign o_code[ 2]   = syndrome_wire[0] ? error_bit[ 6]^x_data_wire[ 2] : x_data_wire[ 2];
        assign o_code[ 1]   = syndrome_wire[0] ? error_bit[ 5]^x_data_wire[ 1] : x_data_wire[ 1];
        assign o_code[ 0]   = syndrome_wire[0] ? error_bit[ 3]^x_data_wire[ 0] : x_data_wire[ 0];
	assign o_parity[7]  = syndrome_wire[0] ? error_bit[64]^x_parity_wire[7]: x_parity_wire[7];
	assign o_parity[6]  = syndrome_wire[0] ? error_bit[32]^x_parity_wire[6]: x_parity_wire[6];
        assign o_parity[5]  = syndrome_wire[0] ? error_bit[16]^x_parity_wire[5]: x_parity_wire[5];
        assign o_parity[4]  = syndrome_wire[0] ? error_bit[8]^x_parity_wire[4]: x_parity_wire[4];
        assign o_parity[3]  = syndrome_wire[0] ? error_bit[4]^x_parity_wire[3]: x_parity_wire[3];
        assign o_parity[2]  = syndrome_wire[0] ? error_bit[2]^x_parity_wire[2]: x_parity_wire[2];
        assign o_parity[1]  = syndrome_wire[0] ? error_bit[1]^x_parity_wire[1]: x_parity_wire[1];
        assign o_parity[0]  = syndrome_wire[0] ? error_bit[0]^x_parity_wire[0]: x_parity_wire[0];	

endmodule

//---------------------------------------------------------------------
// error_bit_decoder module
//---------------------------------------------------------------------
module error_bit_decoder(
    i_data,
    o_decodes
);
parameter data_width = 5;
localparam decodes_width = 1 << data_width;
input  [data_width-1:0]     i_data;
output [decodes_width-1:0]  o_decodes;

reg    [decodes_width-1:0]  o_decodes;

always @(i_data)
begin
    o_decodes = 0;
    o_decodes[i_data] = 1;
end

endmodule

module ecc_dec_wrap (
	o_code,
	o_parity,
	eccoutsberr,
	eccoutdberr,
	i_data,
	i_parity,
	EMB5K_1_PORTA_REG_OUT,
	DEC_REG_EN,
	ECC_DEC_EN,
	c1r1_aa,
	err_addr,
	read_en,
	c1r1_rstna,
	peek_en,
	FIFO_EN,
	PEEK_MODE,
	peek_rd_en,
	c1r1_reg_ena,
	clkreg_a
);

output	[63:0]	o_code;
output	[7:0]	o_parity;
output		eccoutsberr;
output		eccoutdberr;
input	[63:0]	i_data;
input	[7:0] 	i_parity;
input		EMB5K_1_PORTA_REG_OUT;
input		DEC_REG_EN;
input		ECC_DEC_EN;
input   [11:0]  c1r1_aa;
output  [7:0]   err_addr;
input           read_en;
input           c1r1_rstna;
input           peek_en;
input           FIFO_EN;
input           PEEK_MODE;
input           peek_rd_en;
input           c1r1_reg_ena;
input		clkreg_a;

reg        eccoutdberr_reg0_t0;
reg        eccoutsberr_reg0_t0;
reg        eccoutdberr_reg0_t1;
reg        eccoutsberr_reg0_t1;
reg        read_en_reg0;
reg        read_en_reg1;
wire       read_en_mux = DEC_REG_EN ? read_en_reg1 : read_en_reg0;
wire [7:0] c1r1_aa_t = c1r1_aa[11:4];
reg  [7:0] c1r1_aa_reg0;
reg  [7:0] c1r1_aa_reg1_t0;
reg  [7:0] c1r1_aa_reg2_t0;
reg  [7:0] c1r1_aa_reg1_t1;
reg  [7:0] c1r1_aa_reg2_t1;

ECC_DECODER u0 (
	.i_data		(i_data[63:0]),
	.i_parity	(i_parity[7:0]),

	.eccoutdberr	(eccoutdberr_t),
	.eccoutsberr	(eccoutsberr_t),
	.o_code		(o_code[63:0]),
	.o_parity	(o_parity[7:0]) 
);

wire peek_en_n = !peek_en;
wire peek_rd_en_t = FIFO_EN & PEEK_MODE ? peek_rd_en : 1'b1;

always@(posedge clkreg_a or negedge c1r1_rstna)
begin
    if(~c1r1_rstna)
    begin
        eccoutsberr_reg0_t0 <= 0;
        eccoutdberr_reg0_t0 <= 0;
    end
    else if(c1r1_reg_ena)
    begin
        eccoutsberr_reg0_t0 <= eccoutsberr_t & read_en_mux & ECC_DEC_EN;
        eccoutdberr_reg0_t0 <= eccoutdberr_t & read_en_mux & ECC_DEC_EN;
    end
end

always@(posedge clkreg_a or negedge c1r1_rstna)
begin
    if(~c1r1_rstna)
    begin
        eccoutsberr_reg0_t1 <= 0;
        eccoutdberr_reg0_t1 <= 0;
    end
    else if(peek_en_n)
    begin
        eccoutsberr_reg0_t1 <= eccoutsberr_t & read_en_mux & ECC_DEC_EN;
        eccoutdberr_reg0_t1 <= eccoutdberr_t & read_en_mux & ECC_DEC_EN;
    end
end

always@(posedge clkreg_a or negedge c1r1_rstna)
begin
    if(~c1r1_rstna)
    begin
        c1r1_aa_reg1_t0 <= 0;
        c1r1_aa_reg2_t0 <= 0;
    end
    else if(c1r1_reg_ena)
    begin
        c1r1_aa_reg1_t0 <= c1r1_aa_reg0;
        c1r1_aa_reg2_t0 <= c1r1_aa_reg1_t0;
    end
end

always@(posedge clkreg_a or negedge c1r1_rstna)
begin
    if(~c1r1_rstna)
    begin
        c1r1_aa_reg1_t1 <= 0;
        c1r1_aa_reg2_t1 <= 0;
    end
    else if(peek_en_n)
    begin
        c1r1_aa_reg1_t1 <= c1r1_aa_reg0;
        c1r1_aa_reg2_t1 <= c1r1_aa_reg1_t1;
    end
end

always@(posedge clkreg_a or negedge c1r1_rstna)
begin
    if(~c1r1_rstna)
    begin
        read_en_reg0 <= 0;
        c1r1_aa_reg0 <= 0;
    end
    else if(read_en)
    begin
        read_en_reg0 <= read_en;
        c1r1_aa_reg0 <= c1r1_aa_t;
    end
end

always@(posedge clkreg_a or negedge c1r1_rstna)
begin
    if(~c1r1_rstna)
        read_en_reg1 <= 0;
    else
        read_en_reg1 <= read_en_reg0;
end

assign eccoutdberr = EMB5K_1_PORTA_REG_OUT ? peek_rd_en_t ? eccoutdberr_reg0_t0 : eccoutdberr_reg0_t1
                                           : eccoutdberr_t & read_en_mux & ECC_DEC_EN;

assign eccoutsberr = EMB5K_1_PORTA_REG_OUT ? peek_rd_en_t ? eccoutsberr_reg0_t0 : eccoutsberr_reg0_t1
                                           : eccoutsberr_t & read_en_mux & ECC_DEC_EN;

assign err_addr = EMB5K_1_PORTA_REG_OUT ? DEC_REG_EN ? peek_rd_en_t ? c1r1_aa_reg2_t0 : c1r1_aa_reg2_t1
                                                     : peek_rd_en_t ? c1r1_aa_reg1_t0 : c1r1_aa_reg1_t1
                                        : c1r1_aa_reg0;

endmodule

//================================================================================
// Copyright (c) 2012 Capital-micro, Inc.(Beijing)  All rights reserved.
//
// Capital-micro, Inc.(Beijing) Confidential.
//
// No part of this code may be reproduced, distributed, transmitted,
// transcribed, stored in a retrieval system, or translated into any
// human or computer language, in any form or by any means, electronic,
// mechanical, magnetic, manual, or otherwise, without the express
// written permission of Capital-micro, Inc.
//
//================================================================================
// Module Description: 
// This is the encoder module of the ECC IP 
//================================================================================
// Revision History :
//     V1.0   2012-11-30  FPGA IP Grp, first created
//================================================================================
module ECC_ENCODER(
    din,
    eccindberr,
    eccinsberr,
    dino,
    eccpout,
    ECC_ENC_EN
);

//---------------------------------------------------------------------
// inputs & outputs
//---------------------------------------------------------------------
input   [63:0]  din;
output  [63:0]  dino;
output  [7:0] eccpout;

input eccindberr;
input eccinsberr;

input  ECC_ENC_EN;

wire [63:0] i_data;
assign i_data = {64{ECC_ENC_EN}} & din;

wire [71:0] code_wire;
wire [71:0] o_codes;

assign o_codes    = code_wire;

assign eccpout = {o_codes[64],o_codes[32],o_codes[16],o_codes[8],o_codes[4],o_codes[2],o_codes[1],o_codes[0]};

assign dino[63] = din[63];
assign dino[62] = (eccindberr) ? ~din[62] : din[62];
assign dino[61:31] = din[61:31];
assign dino[30] = (eccinsberr || eccindberr) ? ~din[30] : din[30];
assign dino[29:0] = din[29:0];


//---------------------------------------------------------------------
// instantiate module
//---------------------------------------------------------------------
ecc_encoder_core inst_ecc_encoder_core(
    .i_data(i_data),
    .o_code(code_wire)
);
endmodule


//---------------------------------------------------------------------
// Core ECC encoder module
//---------------------------------------------------------------------
module ecc_encoder_core(
    i_data,
    o_code
);

input   [63:0]  i_data;
output  [71:0]  o_code;

wire [71:0]     x;

assign o_code = x;

        //data
        assign x[71:65] = i_data[63:57];
        assign x[63:33] = i_data[56:26];
        assign x[31:17] = i_data[25:11];
        assign x[15: 9] = i_data[10:4];
        assign x[ 7: 5] = i_data[3:1];
        assign x[ 3]    = i_data[0];
        //parity
        assign x[64]    = ^x[71:65];
        assign x[32]    = ^x[63:33];
        assign x[16]    = (^x[63:48])^(^x[31:17]);
        assign x[ 8]    = (^x[63:56])^(^x[47:40])^(^x[31:24])^(^x[15:9]);
        assign x[ 4]    = (^x[71:68])^(^x[63:60])^(^x[55:52])^(^x[47:44])^(^x[39:36])^(^x[31:28])^(^x[23:20])^(^x[15:12])^(^x[7:5]);
        assign x[ 2]    = (^x[71:70])^(^x[67:66])^(^x[63:62])^(^x[59:58])^(^x[55:54])^(^x[51:50])^(^x[47:46])^(^x[43:42])^(^x[39:38])^(^x[35:34])^(^x[31:30])^(^x[27:26])^(^x[23:22])^(^x[19:18])^(^x[15:14])^(^x[11:10])^(^x[7:6])^x[3];
        assign x[ 1]    = x[71]^x[69]^x[67]^x[65]^x[63]^x[61]^x[59]^x[57]^x[55]^x[53]^x[51]^x[49]^x[47]^x[45]^x[43]^x[41]^x[39]^x[37]^x[35]^x[33]^x[31]^x[29]^x[27]^x[25]^x[23]^x[21]^x[19]^x[17]^x[15]^x[13]^x[11]^x[9]^x[7]^x[5]^x[3];
        //extra-parity-bit
        assign x[ 0]    = ^x[71:1];

endmodule

module ecc_enc_wrap (
	dino,
	dinpo,
	ECC_ENC_EN,
	din,
	dinp,
	eccindberr,
	eccinsberr 
);

output	[63:0]	dino;
output	[7:0]	dinpo;
input		ECC_ENC_EN;
input	[63:0]	din;
input	[7:0] 	dinp;
input		eccindberr;
input		eccinsberr;

wire [7:0] eccpout;

ECC_ENCODER ECC_ENCODER (
	.din		(din[63:0]),
	.eccindberr	(eccindberr),
	.eccinsberr	(eccinsberr),
	.ECC_ENC_EN	(ECC_ENC_EN),

	.dino		(dino[63:0]),
	.eccpout	(eccpout[7:0]) 
);

assign dinpo = ECC_ENC_EN ? eccpout[7:0] : dinp[7:0];

endmodule

module emb18k_ext(
     a_addr_ext
    ,b_addr_ext
    ,c1r1_cea_i
    ,c1r1_wea_i
    ,c1r1_ceb_i
    ,c1r1_web_i
    ,c1r2_cea_i
    ,c1r2_wea_i
    ,c1r2_ceb_i
    ,c1r2_web_i
    ,c1r3_cea_i
    ,c1r3_wea_i
    ,c1r3_ceb_i
    ,c1r3_web_i
    ,c1r4_cea_i
    ,c1r4_wea_i
    ,c1r4_ceb_i
    ,c1r4_web_i
    ,c1r1_cea
    ,c1r1_wea
    ,c1r1_ceb
    ,c1r1_web
    ,c1r2_cea
    ,c1r2_wea
    ,c1r2_ceb
    ,c1r2_web
    ,c1r3_cea
    ,c1r3_wea
    ,c1r3_ceb
    ,c1r3_web
    ,c1r4_cea
    ,c1r4_wea
    ,c1r4_ceb
    ,c1r4_web
    ,c1r1_clka
    ,c1r1_clkb
    ,c1r2_clka
    ,c1r2_clkb
    ,c1r3_clka
    ,c1r3_clkb
    ,c1r4_clka
    ,c1r4_clkb
    ,c1r1_rstna
    ,c1r1_rstnb
    ,c1r2_rstna
    ,c1r2_rstnb
    ,c1r3_rstna
    ,c1r3_rstnb
    ,c1r4_rstna
    ,c1r4_rstnb
    ,c1r1_reg_ena
    ,c1r1_reg_enb
    ,c1r2_reg_ena
    ,c1r2_reg_enb
    ,c1r3_reg_ena
    ,c1r3_reg_enb
    ,c1r4_reg_ena
    ,c1r4_reg_enb
    ,gbl_clear_b
    ,modeax18_1
    ,modebx18_1
    ,modeax18_2
    ,modebx18_2
    ,modeax18_3
    ,modebx18_3
    ,modeax18_4
    ,modebx18_4
    ,EMB5K_1_MODEA_SEL
    ,EMB5K_3_MODEA_SEL
    ,EMB5K_1_PORTA_WR_MODE
    ,EMB5K_1_PORTB_WR_MODE
    ,EMB5K_3_PORTA_WR_MODE
    ,EMB5K_3_PORTB_WR_MODE
    ,WIDTH_EXT_MODE01
    ,WIDTH_EXT_MODE23
    ,DEPTH_EXT_MODE01
    ,DEPTH_EXT_MODE23
    ,FIFO_EN
    ,PEEK_MODE
    ,EXT_18K
    ,EMB5K_1_PORTA_REG_OUT
    ,EMB5K_1_PORTB_REG_OUT
    ,EMB5K_2_PORTA_REG_OUT
    ,EMB5K_2_PORTB_REG_OUT
    ,EMB5K_3_PORTA_REG_OUT
    ,EMB5K_3_PORTB_REG_OUT
    ,EMB5K_4_PORTA_REG_OUT
    ,EMB5K_4_PORTB_REG_OUT
//    ,EMB5K_1_PORTA_CKEN
//    ,EMB5K_1_PORTB_CKEN
//    ,EMB5K_2_PORTA_CKEN
//    ,EMB5K_2_PORTB_CKEN
//    ,EMB5K_3_PORTA_CKEN
//    ,EMB5K_3_PORTB_CKEN
//    ,EMB5K_4_PORTA_CKEN
//    ,EMB5K_4_PORTB_CKEN
    ,rd_mem_n
    ,wr_mem_n
    ,rptr
    ,wptr
    ,peek_rd_en
    ,peek_en
    ,c1r1_aa_i
    ,c1r1_ab_i
    ,c1r2_aa_i
    ,c1r2_ab_i
    ,c1r3_aa_i
    ,c1r3_ab_i
    ,c1r4_aa_i
    ,c1r4_ab_i
    ,c1r1_aa
    ,c1r1_ab
    ,c1r2_aa
    ,c1r2_ab
    ,c1r3_aa
    ,c1r3_ab
    ,c1r4_aa
    ,c1r4_ab
    ,c1r1_da_i
    ,c1r1_db_i
    ,c1r2_da_i
    ,c1r2_db_i
    ,c1r3_da_i
    ,c1r3_db_i
    ,c1r4_da_i
    ,c1r4_db_i
    ,c1r1_da
    ,c1r1_db
    ,c1r2_da
    ,c1r2_db
    ,c1r3_da
    ,c1r3_db
    ,c1r4_da
    ,c1r4_db
    ,c1r1_q_i
    ,c1r2_q_i
    ,c1r3_q_i
    ,c1r4_q_i
    ,c1r1_q
    ,c1r2_q
    ,c1r3_q
    ,c1r4_q
    ,c1r1_no_a
    ,c1r1_rstna_t
);

input  [1:0]     a_addr_ext;
input  [1:0]     b_addr_ext;
input            c1r1_cea_i;
input     	 c1r1_wea_i;
input            c1r1_ceb_i;
input   	 c1r1_web_i;
input            c1r2_cea_i;
input	         c1r2_wea_i;
input            c1r2_ceb_i;
input            c1r2_web_i;
input            c1r3_cea_i;
input            c1r3_wea_i;
input            c1r3_ceb_i;
input            c1r3_web_i;
input            c1r4_cea_i;
input            c1r4_wea_i;
input            c1r4_ceb_i;
input            c1r4_web_i;
input            c1r1_clka;
input            c1r1_clkb;
input            c1r2_clka;
input            c1r2_clkb;
input            c1r3_clka;
input            c1r3_clkb;
input            c1r4_clka;
input            c1r4_clkb;
input            c1r1_rstna;
input            c1r1_rstnb;
input            c1r2_rstna;
input            c1r2_rstnb;
input            c1r3_rstna;
input            c1r3_rstnb;
input            c1r4_rstna;
input            c1r4_rstnb;
input            c1r1_reg_ena;
input            c1r1_reg_enb;
input            c1r2_reg_ena;
input            c1r2_reg_enb;
input            c1r3_reg_ena;
input            c1r3_reg_enb;
input            c1r4_reg_ena;
input            c1r4_reg_enb;
input		 gbl_clear_b;
output           c1r1_cea;
output           c1r1_wea;
output           c1r1_ceb;
output           c1r1_web;
output           c1r2_cea;
output           c1r2_wea;
output           c1r2_ceb;
output           c1r2_web;
output           c1r3_cea;
output           c1r3_wea;
output           c1r3_ceb;
output           c1r3_web;
output           c1r4_cea;
output           c1r4_wea;
output           c1r4_ceb;
output           c1r4_web;
input            modeax18_1;
input            modebx18_1;
input            modeax18_2;
input            modebx18_2;
input            modeax18_3;
input            modebx18_3;
input            modeax18_4;
input            modebx18_4;
input  [3:0]     EMB5K_1_MODEA_SEL;
input  [3:0]     EMB5K_3_MODEA_SEL;
input  [1:0]     EMB5K_1_PORTA_WR_MODE;
input  [1:0]     EMB5K_1_PORTB_WR_MODE;
input  [1:0]     EMB5K_3_PORTA_WR_MODE;
input  [1:0]     EMB5K_3_PORTB_WR_MODE;
input            WIDTH_EXT_MODE01;
input            WIDTH_EXT_MODE23;
input            DEPTH_EXT_MODE01;
input            DEPTH_EXT_MODE23;
input            FIFO_EN;
input		 PEEK_MODE;
input            EXT_18K;
input            EMB5K_1_PORTA_REG_OUT;
input            EMB5K_1_PORTB_REG_OUT;
input            EMB5K_2_PORTA_REG_OUT;
input            EMB5K_2_PORTB_REG_OUT;
input            EMB5K_3_PORTA_REG_OUT;
input            EMB5K_3_PORTB_REG_OUT;
input            EMB5K_4_PORTA_REG_OUT;
input            EMB5K_4_PORTB_REG_OUT;
//input            EMB5K_1_PORTA_CKEN;
//input            EMB5K_1_PORTB_CKEN;
//input            EMB5K_2_PORTA_CKEN;
//input            EMB5K_2_PORTB_CKEN;
//input            EMB5K_3_PORTA_CKEN;
//input            EMB5K_3_PORTB_CKEN;
//input            EMB5K_4_PORTA_CKEN;
//input            EMB5K_4_PORTB_CKEN;
input            rd_mem_n;
input            wr_mem_n;
input 		 peek_en;
input		 peek_rd_en;
input   [13:0]   rptr;
input   [13:0]   wptr;
input   [11:0]   c1r1_aa_i;
input   [11:0]   c1r1_ab_i;
input   [11:0]   c1r2_aa_i;
input   [11:0]   c1r2_ab_i;
input   [11:0]   c1r3_aa_i;
input   [11:0]   c1r3_ab_i;
input   [11:0]   c1r4_aa_i;
input   [11:0]   c1r4_ab_i;
output  [11:0]   c1r1_aa;
output  [11:0]   c1r1_ab;
output  [11:0]   c1r2_aa;
output  [11:0]   c1r2_ab;
output  [11:0]   c1r3_aa;
output  [11:0]   c1r3_ab;
output  [11:0]   c1r4_aa;
output  [11:0]   c1r4_ab;
input   [17:0]   c1r1_da_i;
input   [17:0]   c1r1_db_i;
input   [17:0]   c1r2_da_i;
input   [17:0]   c1r2_db_i;
input   [17:0]   c1r3_da_i;
input   [17:0]   c1r3_db_i;
input   [17:0]   c1r4_da_i;
input   [17:0]   c1r4_db_i;
output  [17:0]   c1r1_da;
output  [17:0]   c1r1_db;
output  [17:0]   c1r2_da;
output  [17:0]   c1r2_db;
output  [17:0]   c1r3_da;
output  [17:0]   c1r3_db;
output  [17:0]   c1r4_da;
output  [17:0]   c1r4_db;
input   [17:0]   c1r1_q_i;
input   [17:0]   c1r2_q_i;
input   [17:0]   c1r3_q_i;
input   [17:0]   c1r4_q_i;
output  [17:0]   c1r1_q;
output  [17:0]   c1r2_q;
output  [17:0]   c1r3_q;
output  [17:0]   c1r4_q;
output           c1r1_no_a;
output           c1r1_rstna_t;

//reg  [17:0] c1r1_q_reg;
//reg  [17:0] c1r2_q_reg;
//reg  [17:0] c1r3_q_reg;
//reg  [17:0] c1r4_q_reg;

wire [1:0]  aa_ext = FIFO_EN ? rptr[13:12] : a_addr_ext;
wire [1:0]  ab_ext = FIFO_EN ? wptr[13:12] : b_addr_ext;

wire [1:0] aa_ext01;
wire [1:0] aa_ext23;
wire [1:0] ab_ext01;
wire [1:0] ab_ext23;

wire cfg_ext01 = DEPTH_EXT_MODE01 || WIDTH_EXT_MODE01;
wire cfg_ext23 = DEPTH_EXT_MODE23 || WIDTH_EXT_MODE23;

// CE
assign aa_ext01[0] = EXT_18K ?  aa_ext[0] : aa_ext[0];
assign aa_ext01[1] = EXT_18K ? ~aa_ext[1] : 1'b1;
assign aa_ext23[0] = EXT_18K ?  aa_ext[0] : a_addr_ext[1];
assign aa_ext23[1] = EXT_18K ?  aa_ext[1] : 1'b1;

wire cas_cea01 = FIFO_EN ? ~rd_mem_n : c1r1_cea_i;
wire cas_cea23 = EXT_18K ? cas_cea01 : c1r3_cea_i;

wire c1r1_cea = DEPTH_EXT_MODE01 ? ~aa_ext01[0] & aa_ext01[1] & cas_cea01
                                 : WIDTH_EXT_MODE01 ? cas_cea01
                                                    : cas_cea01;

wire c1r2_cea = DEPTH_EXT_MODE01 ? aa_ext01[0] & aa_ext01[1] & cas_cea01
                                 : WIDTH_EXT_MODE01 ? cas_cea01
                                                    : c1r2_cea_i;

wire c1r3_cea = DEPTH_EXT_MODE23 ? ~aa_ext23[0] & aa_ext23[1] & cas_cea23
                                 : WIDTH_EXT_MODE23 ? cas_cea23
                                                    : c1r3_cea_i;

wire c1r4_cea = DEPTH_EXT_MODE23 ? aa_ext23[0] & aa_ext23[1] & cas_cea23
                                 : WIDTH_EXT_MODE23 ? cas_cea23
                                                    : c1r4_cea_i;

assign ab_ext01[0] = EXT_18K ?  ab_ext[0] : ab_ext[0];
assign ab_ext01[1] = EXT_18K ? ~ab_ext[1] : 1'b1;
assign ab_ext23[0] = EXT_18K ?  ab_ext[0] : b_addr_ext[1];
assign ab_ext23[1] = EXT_18K ?  ab_ext[1] : 1'b1;

wire cas_ceb01 = FIFO_EN ? ~wr_mem_n : c1r1_ceb_i;
wire cas_ceb23 = EXT_18K ? cas_ceb01 : c1r3_ceb_i;

wire c1r1_ceb = DEPTH_EXT_MODE01 ? ~ab_ext01[0] & ab_ext01[1] & cas_ceb01
                                 : WIDTH_EXT_MODE01 ? cas_ceb01
                                                    : cas_ceb01;

wire c1r2_ceb = DEPTH_EXT_MODE01 ? ab_ext01[0] & ab_ext01[1] & cas_ceb01
                                 : WIDTH_EXT_MODE01 ? cas_ceb01
                                                    : c1r2_ceb_i;

wire c1r3_ceb = DEPTH_EXT_MODE23 ? ~ab_ext23[0] & ab_ext23[1] & cas_ceb23
                                 : WIDTH_EXT_MODE23 ? cas_ceb23
                                                    : c1r3_ceb_i;

wire c1r4_ceb = DEPTH_EXT_MODE23 ? ab_ext23[0] & ab_ext23[1] & cas_ceb23
                                 : WIDTH_EXT_MODE23 ? cas_ceb23
                                                    : c1r4_ceb_i;

// WE
wire  c1r1_wea_t = modeax18_1 ? c1r1_wea_i : c1r1_wea_i;
wire  c1r2_wea_t = modeax18_2 ? c1r2_wea_i : c1r2_wea_i;
wire  c1r3_wea_t = modeax18_3 ? c1r3_wea_i : c1r3_wea_i;
wire  c1r4_wea_t = modeax18_4 ? c1r4_wea_i : c1r4_wea_i;

wire  cas_wea01 = FIFO_EN ? 1'b0      : c1r1_wea_t;
wire  cas_wea23 = EXT_18K ? cas_wea01 : c1r3_wea_t;

wire  c1r1_wea,c1r2_wea,c1r3_wea,c1r4_wea;
assign c1r1_wea = DEPTH_EXT_MODE01 | (WIDTH_EXT_MODE01 & FIFO_EN) ? cas_wea01 : cas_wea01;
assign c1r2_wea = DEPTH_EXT_MODE01 | (WIDTH_EXT_MODE01 & FIFO_EN) ? cas_wea01 : c1r2_wea_t;
assign c1r3_wea = DEPTH_EXT_MODE23 | (WIDTH_EXT_MODE23 & FIFO_EN & EXT_18K) ? cas_wea23 : c1r3_wea_t;
assign c1r4_wea = DEPTH_EXT_MODE23 | (WIDTH_EXT_MODE23 & FIFO_EN & EXT_18K) ? cas_wea23 : c1r4_wea_t;

wire  c1r1_web_t = modebx18_1 ? c1r1_web_i : c1r1_web_i;
wire  c1r2_web_t = modebx18_2 ? c1r2_web_i : c1r2_web_i;
wire  c1r3_web_t = modebx18_3 ? c1r3_web_i : c1r3_web_i;
wire  c1r4_web_t = modebx18_4 ? c1r4_web_i : c1r4_web_i;

wire  cas_web01 = FIFO_EN ? {~wr_mem_n}    : c1r1_web_t;
wire  cas_web23 = EXT_18K ? cas_web01      : c1r3_web_t;

wire  c1r1_web,c1r2_web,c1r3_web,c1r4_web;
assign c1r1_web = DEPTH_EXT_MODE01 | (WIDTH_EXT_MODE01 & FIFO_EN) ? cas_web01 : cas_web01;
assign c1r2_web = DEPTH_EXT_MODE01 | (WIDTH_EXT_MODE01 & FIFO_EN) ? cas_web01 : c1r2_web_t;
assign c1r3_web = DEPTH_EXT_MODE23 | (WIDTH_EXT_MODE23 & FIFO_EN & EXT_18K) ? cas_web23 : c1r3_web_t;
assign c1r4_web = DEPTH_EXT_MODE23 | (WIDTH_EXT_MODE23 & FIFO_EN & EXT_18K) ? cas_web23 : c1r4_web_t;

// addr
wire [11:0] cas_aa01 = FIFO_EN ? rptr[11:0] : c1r1_aa_i;
wire [11:0] cas_aa23 = EXT_18K ? cas_aa01   : c1r3_aa_i;

wire [11:0]   c1r1_aa;
wire [11:0]   c1r2_aa;
wire [11:0]   c1r3_aa;
wire [11:0]   c1r4_aa;

assign c1r1_aa = cfg_ext01 ? cas_aa01 : cas_aa01;
assign c1r2_aa = cfg_ext01 ? cas_aa01 : c1r2_aa_i;
assign c1r3_aa = cfg_ext23 ? cas_aa23 : c1r3_aa_i;
assign c1r4_aa = cfg_ext23 ? cas_aa23 : c1r4_aa_i;

wire [11:0] cas_ab01 = FIFO_EN ? wptr[11:0] : c1r1_ab_i;
wire [11:0] cas_ab23 = EXT_18K ? cas_ab01   : c1r3_ab_i;

wire [11:0]   c1r1_ab;
wire [11:0]   c1r2_ab;
wire [11:0]   c1r3_ab;
wire [11:0]   c1r4_ab;

assign c1r1_ab = cfg_ext01 ? cas_ab01 : cas_ab01;
assign c1r2_ab = cfg_ext01 ? cas_ab01 : c1r2_ab_i;
assign c1r3_ab = cfg_ext23 ? cas_ab23 : c1r3_ab_i;
assign c1r4_ab = cfg_ext23 ? cas_ab23 : c1r4_ab_i;

// DI
wire [17:0] cas_da23 = EXT_18K ? c1r1_da_i  : c1r3_da_i;
wire [17:0] c1r1_da;
wire [17:0] c1r2_da;
wire [17:0] c1r3_da;
wire [17:0] c1r4_da;

assign c1r1_da = DEPTH_EXT_MODE01 ? c1r1_da_i : c1r1_da_i;
assign c1r2_da = DEPTH_EXT_MODE01 ? c1r1_da_i : c1r2_da_i;
assign c1r3_da = DEPTH_EXT_MODE23 ? cas_da23  : c1r3_da_i;
assign c1r4_da = DEPTH_EXT_MODE23 ? cas_da23  : c1r4_da_i;

wire [17:0] cas_db23 = EXT_18K ? c1r1_db_i  : c1r3_db_i;
wire [17:0] c1r1_db;
wire [17:0] c1r2_db;
wire [17:0] c1r3_db;
wire [17:0] c1r4_db;

assign c1r1_db = DEPTH_EXT_MODE01 ? c1r1_db_i : c1r1_db_i;
assign c1r2_db = DEPTH_EXT_MODE01 ? c1r1_db_i : c1r2_db_i;
assign c1r3_db = DEPTH_EXT_MODE23 ? cas_db23  : c1r3_db_i;
assign c1r4_db = DEPTH_EXT_MODE23 ? cas_db23  : c1r4_db_i;

// DO
wire [1:0] ab_ext01_t;
wire [1:0] ab_ext23_t;
assign ab_ext01_t[0] = EMB5K_1_MODEA_SEL==4'b0000 ? aa_ext01[0] : ab_ext01[0];
assign ab_ext01_t[1] = ab_ext01[1];
assign ab_ext23_t[0] = EMB5K_3_MODEA_SEL==4'b0000 ? aa_ext23[0] : ab_ext23[0];
assign ab_ext23_t[1] = EMB5K_1_MODEA_SEL==4'b0000 ? aa_ext23[1] : ab_ext23[1];

wire c1r1_regout_ena = EMB5K_1_PORTA_REG_OUT;
wire c1r1_regout_enb = modeax18_1 ? EMB5K_1_PORTA_REG_OUT : EMB5K_1_PORTB_REG_OUT;
wire c1r1_rstna_t = c1r1_rstna & gbl_clear_b;
wire c1r1_rstnb_t = (modeax18_1 ? c1r1_rstna : c1r1_rstnb) & gbl_clear_b;
wire [17:0] c1r1_q_t;
wire [17:0] c1r1_q_tt;
reg aa_ext01_delay0;
reg ab_ext01_delay0;
//peek_rd_en mux
wire peek_rd_en_t = FIFO_EN & PEEK_MODE ? peek_rd_en : 1'b1;


DNT_emb_ckmux2m8 clkb_mux1(.A(c1r1_clkb),.B(c1r1_clka),.S(modeax18_1),  .Z(c1r1_clkreg_b));
//ext addr delay one cycle
//wire c1r1_no_a = (c1r1_cea_i & !c1r1_wea_i)|(c1r1_cea_i & c1r1_wea_i & (EMB5K_1_PORTA_WR_MODE[0] | EMB5K_1_PORTA_WR_MODE[1]));
//wire c1r1_no_b = (c1r1_ceb_i & !c1r1_web_i)|(c1r1_ceb_i & c1r1_web_i & (EMB5K_1_PORTB_WR_MODE[0] | EMB5K_1_PORTB_WR_MODE[1]));
wire c1r1_no_a = (cas_cea01 & !cas_wea01)|(cas_cea01 & cas_wea01 & (EMB5K_1_PORTA_WR_MODE[0] | EMB5K_1_PORTA_WR_MODE[1]));
wire c1r1_no_b = (cas_ceb01 & !cas_web01)|(cas_ceb01 & cas_web01 & (EMB5K_1_PORTB_WR_MODE[0] | EMB5K_1_PORTB_WR_MODE[1]));
//wire c1r1_no_a = (cas_cea01 & !cas_wea01 & !EMB5K_1_PORTA_REG_OUT) |
//                 (cas_cea01 & !cas_wea01 & EMB5K_1_PORTA_REG_OUT & (c1r1_reg_ena|(FIFO_EN&PEEK_MODE))) |
//                 (cas_cea01 & cas_wea01 & (EMB5K_1_PORTA_WR_MODE[0] | EMB5K_1_PORTA_WR_MODE[1]) & !EMB5K_1_PORTA_REG_OUT) |
//                 (cas_cea01 & cas_wea01 & (EMB5K_1_PORTA_WR_MODE[0] | EMB5K_1_PORTA_WR_MODE[1]) & EMB5K_1_PORTA_REG_OUT & (c1r1_reg_ena|(FIFO_EN&PEEK_MODE)));
//wire c1r1_no_b = (cas_ceb01 & !cas_web01 & !EMB5K_1_PORTB_REG_OUT) | 
//                 (cas_ceb01 & !cas_web01 & EMB5K_1_PORTB_REG_OUT & c1r1_reg_enb) | 
//                 (cas_ceb01 & cas_web01 & (EMB5K_1_PORTB_WR_MODE[0] | EMB5K_1_PORTB_WR_MODE[1]) & !EMB5K_1_PORTB_REG_OUT) | 
//                 (cas_ceb01 & cas_web01 & (EMB5K_1_PORTB_WR_MODE[0] | EMB5K_1_PORTB_WR_MODE[1]) & EMB5K_1_PORTB_REG_OUT & c1r1_reg_enb);

wire aa_ext01_en0 = DEPTH_EXT_MODE01 ? c1r1_no_a : 1'b1;
wire ab_ext01_en0 = DEPTH_EXT_MODE01 ? (EMB5K_1_MODEA_SEL==4'b0000 ? c1r1_no_a : c1r1_no_b) : 1'b1;
always@(posedge c1r1_clka or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
	aa_ext01_delay0 <= 1'b0;
    else if(aa_ext01_en0)
	aa_ext01_delay0 <= aa_ext01[0];
end

always@(posedge c1r1_clkreg_b or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
	ab_ext01_delay0 <= 1'b0;
    else if(ab_ext01_en0)
	ab_ext01_delay0 <= ab_ext01_t[0];
end


assign c1r1_q_t[8:0] = aa_ext01_delay0 & DEPTH_EXT_MODE01 ? c1r2_q_i[8:0] : c1r1_q_i[8:0];
assign c1r1_q_t[17:9] = ab_ext01_delay0 & DEPTH_EXT_MODE01 ? c1r2_q_i[17:9] : c1r1_q_i[17:9];


//gclk_clk_and clka_gating1 ( .ck_i0(EMB5K_1_PORTA_CKEN), .ck_i1(c1r1_clka), .ck_out(c1r1_clkreg_a));
//gclk_clk_and clkb_gating1 ( .ck_i0(EMB5K_1_PORTB_CKEN), .ck_i1(c1r1_clkb), .ck_out(c1r1_clkb_t));
//DNT_emb_ckmux2m8 clkb_mux1(.A(c1r1_clkb),.B(c1r1_clka),.S(modeax18_1),  .Z(c1r1_clkreg_b));
reg [17:0] c1r1_q_reg_t0;
reg [17:0] c1r1_q_reg_t1;
wire [17:0] c1r1_q_reg;

always@(posedge c1r1_clka or negedge c1r1_rstna_t)
begin
    if(~c1r1_rstna_t)
        c1r1_q_reg_t0[8:0] <= 9'b0;
    else if(c1r1_reg_ena)
        c1r1_q_reg_t0[8:0] <= c1r1_q_tt[8:0];
end

wire peek_en_n = !peek_en;

always@(posedge c1r1_clka or negedge c1r1_rstna_t)
begin
    if(~c1r1_rstna_t)
        c1r1_q_reg_t1[8:0] <= 9'b0;
    else if(peek_en_n)
        c1r1_q_reg_t1[8:0] <= c1r1_q_tt[8:0];
end

assign c1r1_q_reg[8:0] = peek_rd_en_t ? c1r1_q_reg_t0[8:0] : c1r1_q_reg_t1[8:0];

always@(posedge c1r1_clkreg_b or negedge c1r1_rstnb_t)
begin
    if(~c1r1_rstnb_t)
        c1r1_q_reg_t0[17:9] <= 9'b0;
    else if(c1r1_reg_enb) 
        c1r1_q_reg_t0[17:9] <= c1r1_q_tt[17:9];
end

always@(posedge c1r1_clkreg_b or negedge c1r1_rstnb_t)
begin
    if(~c1r1_rstnb_t)
        c1r1_q_reg_t1[17:9] <= 9'b0;
    else if(peek_en_n)
        c1r1_q_reg_t1[17:9] <= c1r1_q_tt[17:9];
end

assign c1r1_q_reg[17:9] = peek_rd_en_t ? c1r1_q_reg_t0[17:9] : c1r1_q_reg_t1[17:9];


wire c1r2_regout_ena = EMB5K_2_PORTA_REG_OUT;
wire c1r2_regout_enb = modeax18_2 ? EMB5K_2_PORTA_REG_OUT : EMB5K_2_PORTB_REG_OUT;
wire c1r2_rstna_t = c1r2_rstna & gbl_clear_b;
wire c1r2_rstnb_t = (modeax18_2 ? c1r2_rstna : c1r2_rstnb) & gbl_clear_b;

//gclk_clk_and clka_gating2 ( .ck_i0(EMB5K_2_PORTA_CKEN), .ck_i1(c1r2_clka), .ck_out(c1r2_clkreg_a));
//gclk_clk_and clkb_gating2 ( .ck_i0(EMB5K_2_PORTB_CKEN), .ck_i1(c1r2_clkb), .ck_out(c1r2_clkb_t));
DNT_emb_ckmux2m8 clkb_mux2(.A(c1r2_clkb),.B(c1r2_clka),.S(modeax18_2),  .Z(c1r2_clkreg_b));
reg [17:0] c1r2_q_reg_t0;
reg [17:0] c1r2_q_reg_t1;
wire [17:0] c1r2_q_reg;

always@(posedge c1r2_clka or negedge c1r2_rstna_t)
begin
    if(~c1r2_rstna_t)
        c1r2_q_reg_t0[8:0] <= 9'b0;
    else  if(c1r2_reg_ena)
        c1r2_q_reg_t0[8:0] <= c1r2_q_i[8:0];
end

always@(posedge c1r2_clka or negedge c1r2_rstna_t)
begin
    if(~c1r2_rstna_t)
        c1r2_q_reg_t1[8:0] <= 9'b0;
    else if(peek_en_n)
        c1r2_q_reg_t1[8:0] <= c1r2_q_i[8:0];
end

assign c1r2_q_reg[8:0] = peek_rd_en_t ? c1r2_q_reg_t0[8:0] : c1r2_q_reg_t1[8:0];


always@(posedge c1r2_clkreg_b or negedge c1r2_rstnb_t)
begin
    if(~c1r2_rstnb_t)
        c1r2_q_reg_t0[17:9] <= 9'b0;
    else if(c1r2_reg_enb)
        c1r2_q_reg_t0[17:9] <= c1r2_q_i[17:9];
end

always@(posedge c1r2_clkreg_b or negedge c1r2_rstnb_t)
begin
    if(~c1r2_rstnb_t)
        c1r2_q_reg_t1[17:9] <= 9'b0;
    else if(peek_en_n)
        c1r2_q_reg_t1[17:9] <= c1r2_q_i[17:9];
end

assign c1r2_q_reg[17:9] = peek_rd_en_t ? c1r2_q_reg_t0[17:9] : c1r2_q_reg_t1[17:9];



wire c1r3_regout_ena = EMB5K_3_PORTA_REG_OUT;
wire c1r3_regout_enb = modeax18_3 ? EMB5K_3_PORTA_REG_OUT : EMB5K_3_PORTB_REG_OUT;
wire c1r3_rstna_t = c1r3_rstna & gbl_clear_b;
wire c1r3_rstnb_t = (modeax18_3 ? c1r3_rstna : c1r3_rstnb) & gbl_clear_b;
wire [17:0] c1r3_q_t;
reg aa_ext23_delay0;
reg ab_ext23_delay0;
DNT_emb_ckmux2m8 clkb_mux3(.A(c1r3_clkb),.B(c1r3_clka),.S(modeax18_3),  .Z(c1r3_clkreg_b));
//ext addr delay one cycle
//wire c1r3_no_a = (c1r3_cea_i & !c1r3_wea_i)|(c1r3_cea_i & c1r3_wea_i & (EMB5K_3_PORTA_WR_MODE[0] | EMB5K_3_PORTA_WR_MODE[1]));
//wire c1r3_no_b = (c1r3_ceb_i & !c1r3_web_i)|(c1r3_ceb_i & c1r3_web_i & (EMB5K_3_PORTB_WR_MODE[0] | EMB5K_3_PORTB_WR_MODE[1]));
wire c1r3_no_a = (cas_cea23 & !cas_wea23)|(cas_cea23 & cas_wea23 & (EMB5K_3_PORTA_WR_MODE[0] | EMB5K_3_PORTA_WR_MODE[1]));
wire c1r3_no_b = (cas_ceb23 & !cas_web23)|(cas_ceb23 & cas_web23 & (EMB5K_3_PORTB_WR_MODE[0] | EMB5K_3_PORTB_WR_MODE[1]));
//wire c1r3_no_a = (cas_cea23 & !cas_wea23 & !EMB5K_3_PORTA_REG_OUT) |
//                 (cas_cea23 & !cas_wea23 & EMB5K_3_PORTA_REG_OUT & (c1r3_reg_ena|(FIFO_EN&PEEK_MODE&EXT_18K))) |
//                 (cas_cea23 & cas_wea23 & (EMB5K_3_PORTA_WR_MODE[0] | EMB5K_3_PORTA_WR_MODE[1]) & !EMB5K_3_PORTA_REG_OUT) |
//                 (cas_cea23 & cas_wea23 & (EMB5K_3_PORTA_WR_MODE[0] | EMB5K_3_PORTA_WR_MODE[1]) & EMB5K_3_PORTA_REG_OUT & (c1r3_reg_ena|(FIFO_EN&PEEK_MODE&EXT_18K)));
//wire c1r3_no_b = (cas_ceb23 & !cas_web23 & !EMB5K_3_PORTB_REG_OUT) | 
//                 (cas_ceb23 & !cas_web23 & EMB5K_3_PORTB_REG_OUT & c1r3_reg_enb) | 
//                 (cas_ceb23 & cas_web23 & (EMB5K_3_PORTB_WR_MODE[0] | EMB5K_3_PORTB_WR_MODE[1]) & !EMB5K_3_PORTB_REG_OUT) | 
//                 (cas_ceb23 & cas_web23 & (EMB5K_3_PORTB_WR_MODE[0] | EMB5K_3_PORTB_WR_MODE[1]) & EMB5K_3_PORTB_REG_OUT & c1r3_reg_enb);
wire aa_ext23_en0 = DEPTH_EXT_MODE23 ? c1r3_no_a : 1'b1;
wire ab_ext23_en0 = DEPTH_EXT_MODE23 ? (EMB5K_3_MODEA_SEL==4'b0000 ? c1r3_no_a : c1r3_no_b) : 1'b1;

always@(posedge c1r3_clka or negedge gbl_clear_b)
begin 
    if(~gbl_clear_b)
	aa_ext23_delay0 <= 1'b0;
    else if(aa_ext23_en0)
	aa_ext23_delay0 <= aa_ext23[0];
end

always@(posedge c1r3_clkreg_b or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
	ab_ext23_delay0 <= 1'b0;
    else if(ab_ext23_en0)
	ab_ext23_delay0 <= ab_ext23_t[0];
end


assign c1r3_q_t[8:0] = aa_ext23_delay0 & DEPTH_EXT_MODE23 ? c1r4_q_i[8:0] : c1r3_q_i[8:0];
assign c1r3_q_t[17:9] = ab_ext23_delay0 & DEPTH_EXT_MODE23 ? c1r4_q_i[17:9] : c1r3_q_i[17:9];



//gclk_clk_and clka_gating3 ( .ck_i0(EMB5K_3_PORTA_CKEN), .ck_i1(c1r3_clka), .ck_out(c1r3_clkreg_a));
//gclk_clk_and clkb_gating3 ( .ck_i0(EMB5K_3_PORTB_CKEN), .ck_i1(c1r3_clkb), .ck_out(c1r3_clkb_t));
//DNT_emb_ckmux2m8 clkb_mux3(.A(c1r3_clkb),.B(c1r3_clka),.S(modeax18_3),  .Z(c1r3_clkreg_b));
reg [17:0] c1r3_q_reg_t0;
reg [17:0] c1r3_q_reg_t1;
wire [17:0] c1r3_q_reg;

always@(posedge c1r3_clka or negedge c1r3_rstna_t)
begin
    if(~c1r3_rstna_t)
        c1r3_q_reg_t0[8:0] <= 9'b0;
    else if(c1r3_reg_ena)
        c1r3_q_reg_t0[8:0] <= c1r3_q_t[8:0];
end

always@(posedge c1r3_clka or negedge c1r3_rstna_t)
begin
    if(~c1r3_rstna_t)
        c1r3_q_reg_t1[8:0] <= 9'b0;
    else if(peek_en_n)
        c1r3_q_reg_t1[8:0] <= c1r3_q_t[8:0];
end

assign c1r3_q_reg[8:0] = peek_rd_en_t ? c1r3_q_reg_t0[8:0] : c1r3_q_reg_t1[8:0];

always@(posedge c1r3_clkreg_b or negedge c1r3_rstnb_t)
begin
    if(~c1r3_rstnb_t)
        c1r3_q_reg_t0[17:9] <= 9'b0;
    else if(c1r3_reg_enb)
        c1r3_q_reg_t0[17:9] <= c1r3_q_t[17:9];
end

always@(posedge c1r3_clkreg_b or negedge c1r3_rstnb_t)
begin
    if(~c1r3_rstnb_t)
        c1r3_q_reg_t1[17:9] <= 9'b0;
    else if(peek_en_n)
        c1r3_q_reg_t1[17:9] <= c1r3_q_t[17:9];
end

assign c1r3_q_reg[17:9] = peek_rd_en_t ? c1r3_q_reg_t0[17:9] : c1r3_q_reg_t1[17:9];




wire c1r4_regout_ena = EMB5K_4_PORTA_REG_OUT;
wire c1r4_regout_enb = modeax18_4 ? EMB5K_4_PORTA_REG_OUT : EMB5K_4_PORTB_REG_OUT;
wire c1r4_rstna_t = c1r4_rstna & gbl_clear_b;
wire c1r4_rstnb_t = (modeax18_4 ? c1r4_rstna : c1r4_rstnb) & gbl_clear_b;

//gclk_clk_and clka_gating4 ( .ck_i0(EMB5K_4_PORTA_CKEN), .ck_i1(c1r4_clka), .ck_out(c1r4_clkreg_a));
//gclk_clk_and clkb_gating4 ( .ck_i0(EMB5K_4_PORTB_CKEN), .ck_i1(c1r4_clkb), .ck_out(c1r4_clkb_t));
DNT_emb_ckmux2m8 clkb_mux4(.A(c1r4_clkb),.B(c1r4_clka),.S(modeax18_4),  .Z(c1r4_clkreg_b));

reg [17:0] c1r4_q_reg_t0;
reg [17:0] c1r4_q_reg_t1;
wire [17:0] c1r4_q_reg;

always@(posedge c1r4_clka or negedge c1r4_rstna_t)
begin
    if(~c1r4_rstna_t)
        c1r4_q_reg_t0[8:0] <= 9'b0;
    else if(c1r4_reg_ena)
        c1r4_q_reg_t0[8:0] <= c1r4_q_i[8:0];
end

always@(posedge c1r4_clka or negedge c1r4_rstna_t)
begin
    if(~c1r4_rstna_t)
        c1r4_q_reg_t1[8:0] <= 9'b0;
    else if(peek_en_n)
        c1r4_q_reg_t1[8:0] <= c1r4_q_i[8:0];
end

assign c1r4_q_reg[8:0] = peek_rd_en_t ? c1r4_q_reg_t0[8:0] : c1r4_q_reg_t1[8:0];

always@(posedge c1r4_clkreg_b or negedge c1r4_rstnb_t)
begin
    if(~c1r4_rstnb_t)
        c1r4_q_reg_t0[17:9] <= 9'b0;
    else if(c1r4_reg_enb)
        c1r4_q_reg_t0[17:9] <= c1r4_q_i[17:9];
end


always@(posedge c1r4_clkreg_b or negedge c1r4_rstnb_t)
begin
    if(~c1r4_rstnb_t)
        c1r4_q_reg_t1[17:9] <= 9'b0;
    else if(peek_en_n)
        c1r4_q_reg_t1[17:9] <= c1r4_q_i[17:9];
end

assign c1r4_q_reg[17:9] = peek_rd_en_t ? c1r4_q_reg_t0[17:9] : c1r4_q_reg_t1[17:9];

//wire [17:0] c1r1_q_tt;

assign c1r4_q[8:0] = c1r4_regout_ena ? c1r4_q_reg[8:0] : c1r4_q_i[8:0];
assign c1r3_q[8:0] = c1r3_regout_ena ? c1r3_q_reg[8:0] : c1r3_q_t[8:0];

assign c1r2_q[8:0] = c1r2_regout_ena ? c1r2_q_reg[8:0] : c1r2_q_i[8:0];
assign c1r1_q[8:0] = c1r1_regout_ena ? c1r1_q_reg[8:0] : c1r1_q_tt[8:0];
//18K ext addr delay one or two cycles
//reg aa_ext23_delay_1c;
//reg aa_ext23_delay_2c;
//wire aa_ext23_delay1;
//
//wire aa_ext23_en1 = (EXT_18K & DEPTH_EXT_MODE01 & DEPTH_EXT_MODE23) ? c1r1_no_a : 1'b1;
//always@(posedge c1r1_clka or negedge gbl_clear_b)
//begin
//    if(~gbl_clear_b)
//      	aa_ext23_delay_1c <= 1'b0;
//    else if(aa_ext23_en1)
//        aa_ext23_delay_1c <= aa_ext23[1];
//end
//
////reg enable delay one cycle
//reg aa_ext23_en1_delay;
//always@(posedge c1r1_clka or negedge gbl_clear_b)
//begin
//    if(~gbl_clear_b)
//      	aa_ext23_en1_delay <= 1'b0;
//    else 
//        aa_ext23_en1_delay <= aa_ext23_en1;
//end
//
//
//always@(posedge c1r1_clka or negedge gbl_clear_b)
//begin
//    if(~gbl_clear_b)
//      	aa_ext23_delay_2c <= 1'b0;
//    else if(aa_ext23_en1_delay)
//        aa_ext23_delay_2c <= aa_ext23_delay_1c;
//end
//
//assign aa_ext23_delay1 = c1r1_regout_ena? aa_ext23_delay_2c : aa_ext23_delay_1c;
//assign c1r1_q[8:0] = aa_ext23_delay1 & EXT_18K & DEPTH_EXT_MODE01 ? c1r3_q[8:0] : c1r1_q_tt[8:0]; 


assign c1r4_q[17:9] = c1r4_regout_enb ? c1r4_q_reg[17:9] : c1r4_q_i[17:9];
assign c1r3_q[17:9] = c1r3_regout_enb ? c1r3_q_reg[17:9] : c1r3_q_t[17:9];

assign c1r2_q[17:9] = c1r2_regout_enb ? c1r2_q_reg[17:9] : c1r2_q_i[17:9];
assign c1r1_q[17:9] = c1r1_regout_enb ? c1r1_q_reg[17:9] : c1r1_q_tt[17:9];
//18K ext addr delay one or two cycles
//reg ab_ext23_delay_1c;
//reg ab_ext23_delay_2c;
//wire ab_ext23_delay1;
//wire ab_ext23_en1 = (EXT_18K & DEPTH_EXT_MODE01 & DEPTH_EXT_MODE23) ? (EMB5K_1_MODEA_SEL == 4'b0000 ? c1r1_no_a : c1r1_no_b) : 1'b1;
//always@(posedge c1r1_clkreg_b or negedge gbl_clear_b)
//begin
//    if(~gbl_clear_b)
//      	ab_ext23_delay_1c <= 1'b0;
//    else if(ab_ext23_en1)
//        ab_ext23_delay_1c <= ab_ext23_t[1];
//end
//
//
////reg enable delay one cycle
//reg ab_ext23_en1_delay;
//always@(posedge c1r1_clkreg_b or negedge gbl_clear_b)
//begin
//    if(~gbl_clear_b)
//      	ab_ext23_en1_delay <= 1'b0;
//    else 
//        ab_ext23_en1_delay <= ab_ext23_en1;
//end
//
//
//always@(posedge c1r1_clkreg_b or negedge gbl_clear_b)
//begin
//    if(~gbl_clear_b)
//      	ab_ext23_delay_2c <= 1'b0;
//    else if(ab_ext23_en1_delay)
//        ab_ext23_delay_2c <= ab_ext23_delay_1c;
//end
//
//assign ab_ext23_delay1 = c1r1_regout_enb? ab_ext23_delay_2c : ab_ext23_delay_1c;
//assign c1r1_q[17:9] = ab_ext23_delay1 & EXT_18K & DEPTH_EXT_MODE01 ? c1r3_q[17:9] : c1r1_q_tt[17:9]; 

reg aa_ext0123_delay0;
reg ab_ext0123_delay0;

always@(posedge c1r1_clka or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
	aa_ext0123_delay0 <= 1'b0;
    else if(aa_ext01_en0)
	aa_ext0123_delay0 <= aa_ext23[1];
end

always@(posedge c1r1_clkreg_b or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
	ab_ext0123_delay0 <= 1'b0;
    else if(ab_ext01_en0)
	ab_ext0123_delay0 <= ab_ext23_t[1];
end

assign c1r1_q_tt[8:0]  = aa_ext0123_delay0 & EXT_18K ? c1r3_q_t[8:0]  : c1r1_q_t[8:0];
assign c1r1_q_tt[17:9] = ab_ext0123_delay0 & EXT_18K ? c1r3_q_t[17:9] : c1r1_q_t[17:9];


//assign c1r4_q[8:0]  = c1r4_q_i[8:0];
//assign c1r3_q[8:0]  = aa_ext23[0] & DEPTH_EXT_MODE23 ? c1r4_q_i[8:0]
//                                                     : c1r3_q_i[8:0];
//assign c1r2_q[8:0]  = c1r2_q_i[8:0];
//assign c1r1_q[8:0]  = aa_ext23[1] & EXT_18K ? c1r3_q[8:0] 
//                                            : aa_ext01[0] & DEPTH_EXT_MODE01 ? c1r2_q_i[8:0]
//                                                                             : c1r1_q_i[8:0];
//assign c1r4_q[17:9] = c1r4_q_i[17:9];
//assign c1r3_q[17:9] = ab_ext23_t[0] & DEPTH_EXT_MODE23 ? c1r4_q_i[17:9]
//                                                       : c1r3_q_i[17:9];
//assign c1r2_q[17:9] = c1r2_q_i[17:9];
//assign c1r1_q[17:9] = ab_ext23_t[1] & EXT_18K ? c1r3_q[17:9]
//                                              : ab_ext01_t[0] & DEPTH_EXT_MODE01 ? c1r2_q_i[17:9]
//                                                                                 : c1r1_q_i[17:9];

endmodule


module emb5k_core(
     clka
    ,aa
    ,da
    ,cea
    ,wea
    ,clkb
    ,ab
    ,db
    ,ceb
    ,web
    ,q
    ,init_q
    ,MODEA_SEL
    ,MODEB_SEL
    ,PORTA_WR_MODE
    ,PORTB_WR_MODE
    ,DEC_REG_EN
//    ,PORTA_REG_OUT
//    ,PORTB_REG_OUT
    ,PORTA_BYPASS
    ,PORTB_BYPASS
    ,PORTA_CE
    ,PORTB_CE
//    ,PORTA_WE
//    ,PORTB_WE
    ,PORTA_PROG
    ,PORTB_PROG
//    ,PORTA_CKEN
//    ,PORTB_CKEN
    ,modeax18
    ,modebx18
    ,gbl_clear_b
    ,cf_clk
    ,ch1en
    ,initial_en
    ,initial_in
    ,clkreg_a
    ,por_a
    ,por_b
    ,o_code
    ,o_parity
    ,i_data
    ,i_parity
    ,ECC_DEC_EN
);

input          clka;
input  [11:0]  aa;
input  [17:0]  da;
input          cea;
input          wea;
input          clkb;
input  [11:0]  ab;
input  [17:0]  db;
input          ceb;
input          web;
output [17:0]  q;
output [17:0]  init_q;
input  [3:0]   MODEA_SEL;
input  [3:0]   MODEB_SEL;
input  [1:0]   PORTA_WR_MODE;
input  [1:0]   PORTB_WR_MODE;
input          DEC_REG_EN;
//input          PORTA_REG_OUT;
//input          PORTB_REG_OUT;
input	       PORTA_BYPASS;
input	       PORTB_BYPASS;	
input          PORTA_CE;
input          PORTB_CE;
//input          PORTA_WE;
//input          PORTB_WE;
input  [7:0]   PORTA_PROG;
input  [7:0]   PORTB_PROG;
//input          PORTA_CKEN;
//input          PORTB_CKEN;
output         modeax18;
output         modebx18;
input          gbl_clear_b;
input          cf_clk;
input          ch1en;
input          initial_en;
input  [27:0]  initial_in;
output         clkreg_a;
input          por_a;
input	       por_b;
input   [15:0] o_code;
input   [1:0]  o_parity;
output  [15:0] i_data;
output  [1:0]  i_parity;
input          ECC_DEC_EN;

wire  [17:0]   do_b;
wire  [17:0]   do_a;
reg   [17:0]   ox_do;
wire  [17:0]   ox_do_ecc;
wire  [5:0]    cfg_a;
wire  [5:0]    cfg_b;
wire           modeax18;
wire           modebx18;
wire  [3:0]    modeb_s;

wire  [8:0]    wide_9_a;
wire  [8:0]    wide_9_b;
wire  [3:0]    wide_4_a;
wire  [3:0]    wide_4_b;
wire  [1:0]    wide_2_a;
wire  [1:0]    wide_2_b;
wire           wide_1_a;
wire           wide_1_b;
//reg   [17:0]   ox_reg;
wire  [17:0]   q;
wire  [17:0]   init_q;

wire   [11:0]  aa_t;
wire   [17:0]  da_t;
wire           clkreg_a;
wire           clkreg_b;

wire cea_t0 = gbl_clear_b & PORTA_CE & cea;
wire ceb_t0 = gbl_clear_b & PORTB_CE & ceb;
wire wea_t0 = wea;
wire web_t0 = web;

wire cea_t1 = ch1en ? 1'b0 : (initial_en ? initial_in[0] : cea_t0);
wire ceb_t1 = ch1en ? 1'b0 : (initial_en ? 1'b0 : ceb_t0);//when initial, emb5k is sigle port ram.B port dont work
wire wea_t1 = initial_en ? initial_in[1] : wea_t0;
wire web_t1 = web_t0;

assign aa_t = initial_en ? {initial_in[9:2],4'b0000} : aa;
assign da_t = initial_en ? initial_in[27:10] : da;

emb5k_top emb5k_top(
     .ck_a         (clkreg_a)
    ,.ad_a         (aa_t)
    ,.di_a         (da_t)
    ,.ce_a         (cea_t1)
    ,.we_a         (wea_t1)
    ,.cfg_a        ({PORTA_BYPASS,cfg_a})
    ,.do_a         (do_a)
    ,.ck_b         (clkb)
    ,.ad_b         (ab)
    ,.di_b         (db)
    ,.ce_b         (ceb_t1)
    ,.we_b         (web_t1)
    ,.cfg_b        ({PORTB_BYPASS,cfg_b})
    ,.do_b         (do_b)
    ,.papgrm4dmybl (PORTA_PROG)
    ,.pbpgrm4dmybl (PORTB_PROG)
    ,.por_a        (por_a)
    ,.por_b        (por_b)
);

assign wide_9_a = {do_a[17]|do_a[16],do_a[15]|do_a[7],
                    do_a[14]|do_a[6] ,do_a[13]|do_a[5] ,do_a[12]|do_a[4],
                    do_a[11]|do_a[3] ,do_a[10]|do_a[2] ,do_a[9]|do_a[1] ,
                    do_a[8]|do_a[0]};
assign wide_9_b = {do_b[17]|do_b[16],do_b[15]|do_b[7],
                    do_b[14]|do_b[6] ,do_b[13]|do_b[5] ,do_b[12]|do_b[4],
                    do_b[11]|do_b[3] ,do_b[10]|do_b[2] ,do_b[9]|do_b[1] ,
                    do_b[8]|do_b[0]};
assign wide_4_a = {do_a[15]|do_a[11]|do_a[7]|do_a[3],
                   do_a[14]|do_a[10]|do_a[6]|do_a[2],
                   do_a[13]|do_a[9]|do_a[5]|do_a[1],
                   do_a[12]|do_a[8]|do_a[4]|do_a[0]};
assign wide_4_b = {do_b[15]|do_b[11]|do_b[7]|do_b[3],
                   do_b[14]|do_b[10]|do_b[6]|do_b[2],
                   do_b[13]|do_b[9]|do_b[5]|do_b[1],
                   do_b[12]|do_b[8]|do_b[4]|do_b[0]};
assign wide_2_a = {do_a[15]|do_a[13]|do_a[11]|do_a[9]|do_a[7]|do_a[5]|do_a[3]|do_a[1],
                   do_a[14]|do_a[12]|do_a[10]|do_a[8]|do_a[6]|do_a[4]|do_a[2]|do_a[0]};
assign wide_2_b = {do_b[15]|do_b[13]|do_b[11]|do_b[9]|do_b[7]|do_b[5]|do_b[3]|do_b[1],
                   do_b[14]|do_b[12]|do_b[10]|do_b[8]|do_b[6]|do_b[4]|do_b[2]|do_b[0]};

assign wide_1_a ={|do_a[15:0]};
assign wide_1_b ={|do_b[15:0]};

always@(*)
begin
    if(initial_en == 1'b1)
	ox_do[8:0] = do_a[8:0];
    else if({initial_en,MODEA_SEL[3:0]} == 6'b00000)
	ox_do[8:0] = do_a[8:0];
    else if({initial_en,MODEA_SEL[3:0]} == 6'b01000)
	ox_do[8:0] = wide_9_a;
    else if({initial_en,MODEA_SEL[3:0]} == 6'b01100)
	ox_do[8:0] = {5'b0,wide_4_a};
    else if({initial_en,MODEA_SEL[3:0]} == 6'b01110)
	ox_do[8:0] = {7'b0,wide_2_a};
    else if({initial_en,MODEA_SEL[3:0]} == 6'b01111)
	ox_do[8:0] = {8'b0,wide_1_a};
    else
	ox_do[8:0] = wide_9_a;
end

assign modeax18 = MODEA_SEL[3:0]==4'b0000;
assign modebx18 = MODEB_SEL[3:0]==4'b0000;
assign modeb_s[3:0]=modeax18 ? MODEA_SEL[3:0]:MODEB_SEL[3:0];

always@(*)
begin
    if(initial_en == 1'b1)
	ox_do[17:9] = do_a[17:9];
    else if({initial_en,modeb_s[3:0]} == 6'b00000)
	ox_do[17:9] = do_a[17:9];
    else if({initial_en,modeb_s[3:0]} == 6'b01000)
	ox_do[17:9] = wide_9_b;
    else if({initial_en,modeb_s[3:0]} == 6'b01100)
	ox_do[17:9] = {5'b0,wide_4_b};
    else if({initial_en,modeb_s[3:0]} == 6'b01110)
	ox_do[17:9] = {7'b0,wide_2_b};
    else if({initial_en,modeb_s[3:0]} == 6'b01111)
	ox_do[17:9] = {8'b0,wide_1_b};
    else
	ox_do[17:9] = wide_9_b;

end


assign cfg_a = initial_en ? 6'b00_0000 : {PORTA_WR_MODE[1:0],MODEA_SEL[3:0]};
assign cfg_b = initial_en ? 6'b00_0000 : {PORTB_WR_MODE[1:0],MODEB_SEL[3:0]};

//assign regout_ena = PORTA_REG_OUT;
//assign regout_enb = modeax18 ? PORTA_REG_OUT : PORTB_REG_OUT;

//gclk_clk_and clka_gating ( .ck_i0(PORTA_CKEN), .ck_i1(clka), .ck_out(clka_t));
//gclk_clk_and clkb_gating ( .ck_i0(PORTB_CKEN), .ck_i1(clkb), .ck_out(clkb_t));
DNT_emb_ckmux2m8 clka_mux(.A(clka),.B(cf_clk),.S(initial_en),.Z(clkreg_a));
//DNT_emb_ckmux2m8 clkb_mux(.A(clkb),.B(clka),.S(modeax18),  .Z(clkreg_b));

//assign rstna_t = rstna & gbl_clear_b;
//assign rstnb_t = (modeax18 ? rstna : rstnb) & gbl_clear_b;

assign ox_do_ecc = ECC_DEC_EN ? {o_parity[1:0], o_code[15:0]} : ox_do[17:0];

reg  [15:0] i_data_reg;
wire [15:0] i_data_t;
reg  [1:0]  i_parity_reg;
wire [1:0]  i_parity_t;

assign i_data_t   = ECC_DEC_EN ? do_a[15:0]  : 0;
assign i_parity_t = ECC_DEC_EN ? do_a[17:16] : 0;

//DEC_REG_EN;
always@(posedge clkreg_a or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        i_data_reg  <= 0;
    else
        i_data_reg <= i_data_t;
end

always@(posedge clkreg_a or negedge gbl_clear_b)
begin
    if(~gbl_clear_b)
        i_parity_reg  <= 0;
    else
        i_parity_reg <= i_parity_t;
end

assign i_data   = DEC_REG_EN ? i_data_reg   : i_data_t;
assign i_parity = DEC_REG_EN ? i_parity_reg : i_parity_t;

//always@(posedge clkreg_a or negedge rstna_t)
//begin
//    if(~rstna_t)
//        ox_reg[8:0] <= 9'b0;
//    else
//        ox_reg[8:0] <= ox_do_ecc[8:0];
//end
//
//always@(posedge clkreg_b or negedge rstnb_t)
//begin
//    if(~rstnb_t)
//        ox_reg[17:9] <= 9'b0;
//    else
//        ox_reg[17:9] <= ox_do_ecc[17:9];
//end

//assign q[8:0] = initial_en ? ox_do_ecc[8:0] :
//                regout_ena ? ox_reg[8:0]   :
//                             ox_do_ecc[8:0];
//
//assign q[17:9] = initial_en ? ox_do_ecc[17:9] :
//                 regout_enb ? ox_reg[17:9]   :
//                              ox_do_ecc[17:9];

assign q[8:0] = ox_do_ecc[8:0];
assign q[17:9] = ox_do_ecc[17:9];
assign init_q[8:0] = ox_do[8:0];
assign init_q[17:9] = ox_do[17:9];
endmodule

`define HALF_PERIOD
`timescale 1ns/1ns
module emb5k_top(
 ck_a
,ad_a
,di_a
,ce_a
,we_a
,cfg_a
,do_a
,ck_b
,ad_b
,di_b
,ce_b
,we_b
,cfg_b
,do_b
 
,papgrm4dmybl
,pbpgrm4dmybl
,por_a
,por_b
);

input       ck_a;
input [11:0]ad_a;
input [17:0]di_a;
input       ce_a;
input       we_a;
//input [5:0] cfg_a;
input [6:0] cfg_a;	// March 11, 2014 .  Hao added cfg_a[6] for bypass mode
 
input       ck_b;
input [11:0]ad_b;
input [17:0]di_b;
input       ce_b;
input       we_b;
//input [5:0] cfg_b;
input [6:0] cfg_b;	// March 11, 2014 .  Hao added cfg_b[6] for bypass mode
 
output [17:0]do_a;
output [17:0]do_b;
 
input [7:0]papgrm4dmybl;
input [7:0]pbpgrm4dmybl;
input por_a;
input por_b;

reg [17:0] do_a,do_b;
reg [17:0] do_a_comb,do_b_comb;
reg [17:0] do_a_tmp,do_b_tmp;
reg [17:0] di_a_reg,di_b_reg;
reg [11:0] ad_a_reg,ad_b_reg;
reg        ce_a_reg,we_a_reg;
reg        ce_b_reg,we_b_reg;
reg [17:0] tmp_a,tmp_b;
reg [17:0] mem [0:255];
reg [17:0] do_a_first_read;
reg [17:0] do_b_first_read;

wire [11:4] ad_a_reg_tmp;
wire [11:4] ad_b_reg_tmp;
wire bypen_a ;
wire bypen_b ;

// Hao added cfg_a/b[6] for bypass mode on 03/11/2014

assign bypen_a =(ce_a_reg && !we_a_reg && ce_b_reg && we_b_reg && (ad_a_reg[11:4]==ad_b_reg[11:4])) && cfg_a[6];
assign bypen_b =(ce_b_reg && !we_b_reg && ce_a_reg && we_a_reg && (ad_a_reg[11:4]==ad_b_reg[11:4])) && cfg_b[6];
//assign bypen_a =(ce_a_reg && !we_a_reg && ce_b_reg && we_b_reg && (ad_a_reg[11:4]==ad_b_reg[11:4]));
//assign bypen_b =(ce_b_reg && !we_b_reg && ce_a_reg && we_a_reg && (ad_a_reg[11:4]==ad_b_reg[11:4]));
//for read first
always@(posedge ck_a)begin
do_a_first_read<=mem[ad_a[11:4]];
end

always@(posedge ck_b)begin
do_b_first_read<=mem[ad_b[11:4]];
end

//interface registers
always@(negedge por_a or posedge ck_a)begin
if (~por_a)  begin
  ce_a_reg <=1'b0;
  we_a_reg <=1'b0;
  ad_a_reg[11:4] <=8'b0;
  //do_a=do_a;  // Look into it later
end else begin
  ad_a_reg[11:4]<=ad_a[11:4];
  ce_a_reg<=ce_a;
  we_a_reg<=we_a;
end
end

always @(posedge ck_a) begin
  ad_a_reg[3:0] <= ad_a[3:0];
  di_a_reg <= di_a;
end


always@(negedge por_b or posedge ck_b) begin
if (~por_b) begin
  ad_b_reg[11:4] <= 8'b0;
  ce_b_reg <= 1'b0;
  we_b_reg <= 1'b0;
end else begin
  ad_b_reg[11:4]<=ad_b[11:4];
  ce_b_reg<=ce_b;
  we_b_reg<=we_b;
end
end

always @(posedge ck_b) begin
  ad_b_reg[3:0] <= ad_b[3:0];
  di_b_reg <= di_b;
end

assign ad_a_reg_tmp=ad_a_reg[11:4];
assign ad_b_reg_tmp=ad_b_reg[11:4];

//prepare write in data
always@(*)
begin
tmp_a = mem[ad_a_reg_tmp];
if(cfg_a[3:0] == 4'b1111)
begin
       if(ad_a_reg[3:0] == 00)  tmp_a[00] = di_a_reg[00];
  else if(ad_a_reg[3:0] == 01)  tmp_a[01] = di_a_reg[01];
  else if(ad_a_reg[3:0] == 02)  tmp_a[02] = di_a_reg[02];
  else if(ad_a_reg[3:0] == 03)  tmp_a[03] = di_a_reg[03];
  else if(ad_a_reg[3:0] == 04)  begin
  tmp_a[04] = di_a_reg[04];
  tmp_a[16] = di_a_reg[16];
  end
  //else if(ad_a_reg[3:0] == 04)  tmp_a[04] = di_a_reg[04];
  else if(ad_a_reg[3:0] == 04)  tmp_a[04] = di_a_reg[04];
  else if(ad_a_reg[3:0] == 05)  tmp_a[05] = di_a_reg[05];
  else if(ad_a_reg[3:0] == 06)  tmp_a[06] = di_a_reg[06];
  else if(ad_a_reg[3:0] == 07)  tmp_a[07] = di_a_reg[07];
  else if(ad_a_reg[3:0] == 08)  tmp_a[08] = di_a_reg[08];
  else if(ad_a_reg[3:0] == 09)  tmp_a[09] = di_a_reg[09];
  else if(ad_a_reg[3:0] == 10)  tmp_a[10] = di_a_reg[10];
  else if(ad_a_reg[3:0] == 11)  tmp_a[11] = di_a_reg[11];
  else if(ad_a_reg[3:0] == 12)  tmp_a[12] = di_a_reg[12];
  else if(ad_a_reg[3:0] == 13)  begin
  tmp_a[13] = di_a_reg[13];
  tmp_a[17] = di_a_reg[17];
  end
  //else if(ad_a_reg[3:0] == 13)  tmp_a[13] = di_a_reg[13];
  else if(ad_a_reg[3:0] == 14)  tmp_a[14] = di_a_reg[14];
  else                          tmp_a[15] = di_a_reg[15];
end
else if(cfg_a[3:0] == 4'b1110)
begin
       if(ad_a_reg[3:1] == 0)  tmp_a[01:00] = di_a_reg[01:00];
  else if(ad_a_reg[3:1] == 1)  tmp_a[03:02] = di_a_reg[03:02];
  else if(ad_a_reg[3:1] == 2)  begin
  tmp_a[05:04] = di_a_reg[05:04];
  tmp_a[16] = di_a_reg[16];
  end
  //else if(ad_a_reg[3:1] == 2)  tmp_a[05:04] = di_a_reg[05:04];
  else if(ad_a_reg[3:1] == 3)  tmp_a[07:06] = di_a_reg[07:06];
  else if(ad_a_reg[3:1] == 4)  tmp_a[09:08] = di_a_reg[09:08];
  else if(ad_a_reg[3:1] == 5)  tmp_a[11:10] = di_a_reg[11:10];
  else if(ad_a_reg[3:1] == 6)  begin
  tmp_a[13:12] = di_a_reg[13:12];
  tmp_a[17] = di_a_reg[17];
  end
  //else if(ad_a_reg[3:1] == 6)  tmp_a[13:12] = di_a_reg[13:12];
  else                         tmp_a[15:14] = di_a_reg[15:14];
end
else if(cfg_a[3:0] == 4'b1100)
 begin
       if(ad_a_reg[3:2] == 0) tmp_a[03:00] = di_a_reg[03:00];
  else if(ad_a_reg[3:2] == 1) begin
  tmp_a[07:04] = di_a_reg[07:04];
  tmp_a[16] = di_a_reg[16];
  end
  //else if(ad_a_reg[3:2] == 1) tmp_a[07:04] = di_a_reg[07:04];
  else if(ad_a_reg[3:2] == 2) tmp_a[11:08] = di_a_reg[11:08];
  else begin
  tmp_a[15:12] = di_a_reg[15:12];
  tmp_a[17] = di_a_reg[17];
  end
  //else                        tmp_a[15:12] = di_a_reg[15:12];
 end
else if(cfg_a[3:0] == 4'b1000)
 begin
        if(ad_a_reg[3])  {tmp_a[17],tmp_a[15:08]} = {di_a_reg[17],di_a_reg[15:08]};
        else             {tmp_a[16],tmp_a[07:00]} = {di_a_reg[16],di_a_reg[07:00]};
 end
else if(cfg_a[3:0] == 4'b0000)
 tmp_a = di_a_reg;
end

always@(*)
begin
tmp_b = mem[ad_b_reg_tmp];
if(cfg_b[3:0] == 4'b1111)
begin
       if(ad_b_reg[3:0] == 00)  tmp_b[00] = di_b_reg[00];
  else if(ad_b_reg[3:0] == 01)  tmp_b[01] = di_b_reg[01];
  else if(ad_b_reg[3:0] == 02)  tmp_b[02] = di_b_reg[02];
  else if(ad_b_reg[3:0] == 03)  tmp_b[03] = di_b_reg[03];
  else if(ad_b_reg[3:0] == 04)  begin
  tmp_b[04] = di_b_reg[04];
  tmp_b[16] = di_b_reg[16];
  end
  //else if(ad_b_reg[3:0] == 04)  tmp_b[04] = di_b_reg[04];
  else if(ad_b_reg[3:0] == 05)  tmp_b[05] = di_b_reg[05];
  else if(ad_b_reg[3:0] == 06)  tmp_b[06] = di_b_reg[06];
  else if(ad_b_reg[3:0] == 07)  tmp_b[07] = di_b_reg[07];
  else if(ad_b_reg[3:0] == 08)  tmp_b[08] = di_b_reg[08];
  else if(ad_b_reg[3:0] == 09)  tmp_b[09] = di_b_reg[09];
  else if(ad_b_reg[3:0] == 10)  tmp_b[10] = di_b_reg[10];
  else if(ad_b_reg[3:0] == 11)  tmp_b[11] = di_b_reg[11];
  else if(ad_b_reg[3:0] == 12)  tmp_b[12] = di_b_reg[12];
  else if(ad_b_reg[3:0] == 13)  begin
  tmp_b[13] = di_b_reg[13];
  tmp_b[17] = di_b_reg[17];
  end
  //else if(ad_b_reg[3:0] == 13)  tmp_b[13] = di_b_reg[13];
  else if(ad_b_reg[3:0] == 14)  tmp_b[14] = di_b_reg[14];
  else                          tmp_b[15] = di_b_reg[15];
end
else if(cfg_b[3:0] == 4'b1110)
begin
       if(ad_b_reg[3:1] == 0)  tmp_b[01:00] = di_b_reg[01:00];
  else if(ad_b_reg[3:1] == 1)  tmp_b[03:02] = di_b_reg[03:02];
  else if(ad_b_reg[3:1] == 2)  begin
  tmp_b[05:04] = di_b_reg[05:04];
  tmp_b[16] = di_b_reg[16];
  end
  //else if(ad_b_reg[3:1] == 2)  tmp_b[05:04] = di_b_reg[05:04];
  else if(ad_b_reg[3:1] == 3)  tmp_b[07:06] = di_b_reg[07:06];
  else if(ad_b_reg[3:1] == 4)  tmp_b[09:08] = di_b_reg[09:08];
  else if(ad_b_reg[3:1] == 5)  tmp_b[11:10] = di_b_reg[11:10];
  else if(ad_b_reg[3:1] == 6)  begin
  tmp_b[13:12] = di_b_reg[13:12];
  tmp_b[17] = di_b_reg[17];
  end
  //else if(ad_b_reg[3:1] == 6)  tmp_b[13:12] = di_b_reg[13:12];
  else                         tmp_b[15:14] = di_b_reg[15:14];
end
else if(cfg_b[3:0] == 4'b1100)
 begin
       if(ad_b_reg[3:2] == 0) tmp_b[03:00] = di_b_reg[03:00];
  else if(ad_b_reg[3:2] == 1) begin
  tmp_b[07:04] = di_b_reg[07:04];
  tmp_b[16] = di_b_reg[16];
  end
  //else if(ad_b_reg[3:2] == 1) tmp_b[07:04] = di_b_reg[07:04];
  else if(ad_b_reg[3:2] == 2) tmp_b[11:08] = di_b_reg[11:08];
  else begin
  tmp_b[15:12] = di_b_reg[15:12];
  tmp_b[17] = di_b_reg[17];
  end
  //else                        tmp_b[15:12] = di_b_reg[15:12];
 end
else if(cfg_b[3:0] == 4'b1000)
 begin
        if(ad_b_reg[3])  {tmp_b[17],tmp_b[15:08]} = {di_b_reg[17],di_b_reg[15:08]};
        else             {tmp_b[16],tmp_b[07:00]} = {di_b_reg[16],di_b_reg[07:00]};
 end
else if(cfg_b[3:0] == 4'b0000)
 tmp_b = di_b_reg;
end

//write operation  and read operation
always@(*)
begin
 if(ce_a_reg&we_a_reg)//write
   mem[ad_a_reg_tmp]=tmp_a;
end
wire pa_wrf ; // Port a in write first mode
wire pa_rdf ; // Port a in read first mode
wire pb_wrf ; // Port b in write first mode
wire pb_rdf ; // Port b in read first mode

assign pa_wrf = cfg_a[4] & !cfg_a[5] & we_a_reg;
assign pa_rdf = cfg_a[5];
assign pb_wrf = cfg_b[4] & !cfg_b[5] & we_b_reg;
assign pb_rdf = cfg_b[5];

//always@(*)
always@(ce_a_reg or we_a_reg or ad_a_reg_tmp or do_a_first_read or pa_wrf or tmp_a or do_a_tmp)
begin
	if(ce_a_reg)
    // In sdp mode, we_a_reg is always false and we need do_a_first_read to make sure the do_a is previously stored data. 
    // That's why we put the clause "if (cfg_a[5])" before "if (!we_a_reg)".
      if (cfg_a[5]) //read first 
          do_a_tmp = do_a_first_read;
	  else 
	  	if(!we_a_reg)//read
	      do_a_tmp=mem[ad_a_reg_tmp];

	    /*
	    else if (cfg_a[4]) //write through
	    */
	    else if (pa_wrf) //write through
	      do_a_tmp=tmp_a;
	    else do_a_tmp=do_a_tmp;//not write through
	else //no operation
	  do_a_tmp=do_a_tmp;
end

always@(*)
begin
 if(ce_b_reg&we_b_reg)//write
   mem[ad_b_reg_tmp]=tmp_b;
end

//always@(*)
always@(ce_b_reg or we_b_reg or ad_b_reg_tmp or do_b_first_read or pb_wrf or tmp_b or do_b_tmp)
begin
	if(ce_b_reg)
	  if(!we_b_reg)//read
	    do_b_tmp=mem[ad_b_reg_tmp];
	  else //write
      if (cfg_b[5]) //read first
        do_b_tmp= do_b_first_read;
	    /*
	    else if (cfg_b[4])//write through
	    */
	    else if (pb_wrf)//write through
	      do_b_tmp=tmp_b;
	    else do_b_tmp=do_b_tmp;//not write through
	else //no operation
	  do_b_tmp=do_b_tmp;
end

//prepare output data
always@(*)
begin
if(cfg_a[3:0] == 4'b1111)
begin  
    if(ad_a_reg[3:0] == 00)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0000_0001;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_0001;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_0001;
    end
  else if(ad_a_reg[3:0] == 01)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0000_0010;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_0010;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_0010;
      /*
      if(bypen_a) do_a_comb = tmp_b & 18'b00_0000_0000_0000_0010;
      else        do_a_comb = do_a_tmp & 18'b00_0000_0000_0000_0010;
      */
    end
  else if(ad_a_reg[3:0] == 02)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0000_0100;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_0100;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_0100;
      /*
      if(bypen_a) do_a_comb = tmp_b & 18'b00_0000_0000_0000_0100;
      else        do_a_comb = do_a_tmp & 18'b00_0000_0000_0000_0100;
      */
    end
  else if(ad_a_reg[3:0] == 03)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0000_1000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_1000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_1000;
    end
  else if(ad_a_reg[3:0] == 04)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0001_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0001_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0001_0000;
      /*
      if(bypen_a) do_a_comb = tmp_b & 18'b00_0000_0000_0001_0000;
      else        do_a_comb = do_a_tmp & 18'b00_0000_0000_0001_0000;
      */
    end
  else if(ad_a_reg[3:0] == 05)  
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0010_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0010_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0010_0000;
      end
  else if(ad_a_reg[3:0] == 06) 
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0100_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0100_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0100_0000;
    end
  else if(ad_a_reg[3:0] == 07)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_1000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_1000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_1000_0000;
    end
  else if(ad_a_reg[3:0] == 08)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0001_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0001_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0001_0000_0000;
    end
  else if(ad_a_reg[3:0] == 09)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0010_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0010_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0010_0000_0000;
    end
  else if(ad_a_reg[3:0] == 10)  
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0100_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0100_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_0100_0000_0000;
    end
  else if(ad_a_reg[3:0] == 11)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_1000_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_1000_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0000_1000_0000_0000;
    end
  else if(ad_a_reg[3:0] == 12)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0001_0000_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0001_0000_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0001_0000_0000_0000;
    end
  else if(ad_a_reg[3:0] == 13)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0010_0000_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0010_0000_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0010_0000_0000_0000;
    end
  else if(ad_a_reg[3:0] == 14)
    begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_0100_0000_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0100_0000_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_0100_0000_0000_0000;
    end
  else begin
      if(bypen_a) do_a_comb = tmp_b & 18'bxx_1000_0000_0000_0000;
      else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_1000_0000_0000_0000;
      else        do_a_comb = do_a_tmp & 18'bxx_1000_0000_0000_0000;
  end
end
else if(cfg_a[3:0] == 4'b1110) // 2 data width
begin
  if(ad_a_reg[3:1] == 0) 
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0000_0011;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_0011;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_0011;
  end
  else if(ad_a_reg[3:1] == 1) 
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0000_1100;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_1100;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_1100;
    /*
    if(bypen_a) do_a_comb = tmp_b & 18'b00_0000_0000_0000_1100;
    else        do_a_comb = do_a_tmp & 18'b00_0000_0000_0000_1100;
    */
  end
  else if(ad_a_reg[3:1] == 2) 
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_0011_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0011_0000;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_0011_0000;
    /*
    if(bypen_a) do_a_comb = tmp_b & 18'b00_0000_0000_0011_0000;
    else        do_a_comb = do_a_tmp & 18'b00_0000_0000_0011_0000;
    */
  end
  else if(ad_a_reg[3:1] == 3)  
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_1100_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_1100_0000;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_1100_0000;
  end
  else if(ad_a_reg[3:1] == 4) 
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0011_0000_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0011_0000_0000;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_0011_0000_0000;
  end
  else if(ad_a_reg[3:1] == 5)
  begin
    if(bypen_a)  do_a_comb = tmp_b & 18'bxx_0000_1100_0000_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_1100_0000_0000;
    else         do_a_comb = do_a_tmp & 18'bxx_0000_1100_0000_0000;
  end
  else if(ad_a_reg[3:1] == 6)
  begin
    if(bypen_a)  do_a_comb = tmp_b & 18'bxx_0011_0000_0000_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0011_0000_0000_0000;
    else         do_a_comb = do_a_tmp & 18'bxx_0011_0000_0000_0000;
  end
  else begin
    if(bypen_a)  do_a_comb = tmp_b & 18'bxx_1100_0000_0000_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_1100_0000_0000_0000;
    else         do_a_comb = do_a_tmp & 18'bxx_1100_0000_0000_0000;
  end
end
else if(cfg_a[3:0] == 4'b1100)  // 4 bits data width
 begin
  if(ad_a_reg[3:2] == 0)
  begin  
    if(bypen_a)  do_a_comb = tmp_b & 18'bxx_0000_0000_0000_1111;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_0000_1111;
    else         do_a_comb = do_a_tmp & 18'bxx_0000_0000_0000_1111;
  end
  else if(ad_a_reg[3:2] == 1) 
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_0000_1111_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_0000_1111_0000;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_0000_1111_0000;
    //if(bypen_a) do_a_comb = tmp_b & 18'b00_0000_0000_1111_0000;
    //else        do_a_comb = do_a_tmp & 18'b00_0000_0000_1111_0000;
  end
  else if(ad_a_reg[3:2] == 2) 
  begin
    if(bypen_a) do_a_comb = tmp_b & 18'bxx_0000_1111_0000_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_0000_1111_0000_0000;
    else        do_a_comb = do_a_tmp & 18'bxx_0000_1111_0000_0000;
  end
  else begin
    if(bypen_a)      do_a_comb = tmp_b & 18'bxx_1111_0000_0000_0000;
    else if(pa_wrf) do_a_comb = di_a_reg & 18'bxx_1111_0000_0000_0000;
    else             do_a_comb = do_a_tmp & 18'bxx_1111_0000_0000_0000;
    /*
    if(bypen_a) do_a_comb = tmp_b & 18'b00_1111_0000_0000_0000;
    else        do_a_comb = do_a_tmp & 18'b00_1111_0000_0000_0000;
    */
  end
 end
else if(cfg_a[3:0] == 4'b1000)
 begin
     if(~ad_a_reg[3]) begin
	  if(bypen_a) begin
	  do_a_comb =tmp_b & 18'b01_0000_0000_1111_1111;
	  end
	  else begin
	  do_a_comb = do_a_tmp & 18'b01_0000_0000_1111_1111;
	  end
     end
     if(ad_a_reg[3]) begin
          if(bypen_a) begin
	  do_a_comb =tmp_b & 18'b10_1111_1111_0000_0000;
	  end
	  else begin
	  do_a_comb = do_a_tmp & 18'b10_1111_1111_0000_0000;
          end
     end
 end
else if(cfg_a[3:0] == 4'b0000) begin
  if(bypen_a) begin
  do_a_comb = tmp_b;
  end
  else begin
  do_a_comb = do_a_tmp;
  end
end
end

//a port output
always@(*) begin
  if (ck_a && ce_a_reg && por_a)begin
    if(!we_a_reg) begin //read
      if(cfg_a[3:0]== 4'b1100 || cfg_a[3:0]== 4'b1110 || cfg_a[3:0]== 4'b1111) begin
      do_a={2'bx,do_a_comb[15:0]};
      end
      else begin
      do_a=do_a_comb;
      end
    end
    else begin//write
     /*
      if (cfg_a[4]||cfg_a[5]) begin //write_through or read first
      */
      if (pa_wrf || pa_rdf) begin //write_through or read first
        if(cfg_a[3:0]== 4'b1100 || cfg_a[3:0]== 4'b1110 || cfg_a[3:0]== 4'b1111) begin
        do_a={2'bx,do_a_comb[15:0]};
        end
        else begin
	do_a=do_a_comb;
	end
      end

      else begin // write no-change mode
       do_a=do_a ;
      end
    end
 end
 //else if (~por_a) do_a=0;
end 
	  
always@(*)
begin
if(cfg_b[3:0] == 4'b1111)
begin  
    if(ad_b_reg[3:0] == 00)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0000_0001;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_0001;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_0001;
    end
  else if(ad_b_reg[3:0] == 01)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0000_0010;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_0010;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_0010;
    end
  else if(ad_b_reg[3:0] == 02)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0000_0100;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_0100;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_0100;
    end
  else if(ad_b_reg[3:0] == 03)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0000_1000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_1000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_1000;
    end
  else if(ad_b_reg[3:0] == 04)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0001_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0001_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0001_0000;
    end
  else if(ad_b_reg[3:0] == 05)  
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0010_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0010_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0010_0000;
      end
  else if(ad_b_reg[3:0] == 06) 
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0100_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0100_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0100_0000;
    end
  else if(ad_b_reg[3:0] == 07)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_1000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_1000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_1000_0000;
    end
  else if(ad_b_reg[3:0] == 08)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0001_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0001_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0001_0000_0000;
    end
  else if(ad_b_reg[3:0] == 09)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0010_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0010_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0010_0000_0000;
    end
  else if(ad_b_reg[3:0] == 10)  
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0100_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0100_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_0100_0000_0000;
    end
  else if(ad_b_reg[3:0] == 11)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_1000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_1000_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0000_1000_0000_0000;
    end
  else if(ad_b_reg[3:0] == 12)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0001_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0001_0000_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0001_0000_0000_0000;
    end
  else if(ad_b_reg[3:0] == 13)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0010_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0010_0000_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0010_0000_0000_0000;
    end
  else if(ad_b_reg[3:0] == 14)
    begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_0100_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0100_0000_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_0100_0000_0000_0000;
    end
  else begin
      if(bypen_b) do_b_comb = tmp_a & 18'bxx_1000_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_1000_0000_0000_0000;
      else        do_b_comb = do_b_tmp & 18'bxx_1000_0000_0000_0000;
  end
end
else if(cfg_b[3:0] == 4'b1110)
begin
  if(ad_b_reg[3:1] == 0) 
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0000_0011;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_0011;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_0011;
    /*
    if(bypen_b) do_b_comb = tmp_a & 18'b00_0000_0000_0000_0011;
    else        do_b_comb = do_b_tmp & 18'b00_0000_0000_0000_0011;
    */
  end
  else if(ad_b_reg[3:1] == 1) 
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0000_1100;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_1100;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_1100;
  end
  else if(ad_b_reg[3:1] == 2) 
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_0011_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0011_0000;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_0011_0000;
  end
  else if(ad_b_reg[3:1] == 3)  
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_1100_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_1100_0000;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_1100_0000;
  end
  else if(ad_b_reg[3:1] == 4) 
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0011_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0011_0000_0000;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_0011_0000_0000;
  end
  else if(ad_b_reg[3:1] == 5)
  begin
    if(bypen_b)  do_b_comb = tmp_a & 18'bxx_0000_1100_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_1100_0000_0000;
    else         do_b_comb = do_b_tmp & 18'bxx_0000_1100_0000_0000;
  end
  else if(ad_b_reg[3:1] == 6)
  begin
    if(bypen_b)  do_b_comb = tmp_a & 18'bxx_0011_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0011_0000_0000_0000;
    else         do_b_comb = do_b_tmp & 18'bxx_0011_0000_0000_0000;
  end
  else begin
    if(bypen_b)  do_b_comb = tmp_a & 18'bxx_1100_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_1100_0000_0000_0000;
    else         do_b_comb = do_b_tmp & 18'bxx_1100_0000_0000_0000;
  end
end
else if(cfg_b[3:0] == 4'b1100) // 4 bits data width
 begin
  if(ad_b_reg[3:2] == 0)
  begin  
    if(bypen_b)  do_b_comb = tmp_a & 18'bxx_0000_0000_0000_1111;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_0000_1111;
    else         do_b_comb = do_b_tmp & 18'bxx_0000_0000_0000_1111;
    /*
    if(bypen_b)  do_b_comb = tmp_a & 18'b00_0000_0000_0000_1111;
    else         do_b_comb = do_b_tmp & 18'b00_0000_0000_0000_1111;
    */
  end
  else if(ad_b_reg[3:2] == 1) 
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_0000_1111_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_0000_1111_0000;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_0000_1111_0000;
  end
  else if(ad_b_reg[3:2] == 2) 
  begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_0000_1111_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_0000_1111_0000_0000;
    else        do_b_comb = do_b_tmp & 18'bxx_0000_1111_0000_0000;
  end
  else begin
    if(bypen_b) do_b_comb = tmp_a & 18'bxx_1111_0000_0000_0000;
      else if(pb_wrf) do_b_comb = di_b_reg & 18'bxx_1111_0000_0000_0000;
    else        do_b_comb = do_b_tmp & 18'bxx_1111_0000_0000_0000;
  end
 end
else if(cfg_b[3:0] == 4'b1000)
 begin
     if(~ad_b_reg[3]) begin
	  if(bypen_b) begin
	  do_b_comb =tmp_a & 18'b01_0000_0000_1111_1111;
	  end
	  else begin
	  do_b_comb = do_b_tmp & 18'b01_0000_0000_1111_1111;
	  end
     end
     if(ad_b_reg[3]) begin
          if(bypen_b) begin
	  do_b_comb =tmp_a & 18'b10_1111_1111_0000_0000;
	  end
	  else begin
	  do_b_comb = do_b_tmp & 18'b10_1111_1111_0000_0000;
          end
     end
 end
else if(cfg_b[3:0] == 4'b0000) begin
  if(bypen_b) begin
  do_b_comb = tmp_a;
  end
  else begin
  do_b_comb = do_b_tmp;
  end
end
end

always@(*) begin
  if (ck_b && ce_b_reg && por_b)begin
    if(!we_b_reg) begin //read
      if(cfg_b[3:0]== 4'b1100 || cfg_b[3:0]== 4'b1110 || cfg_b[3:0]== 4'b1111) begin
      do_b={2'bx,do_b_comb[15:0]};
      end
      else begin
      do_b=do_b_comb;
      end
    end
    else begin//write
    /*
      if (cfg_b[4]||cfg_b[5]) begin//write_through or read first
    */
      if ( pb_wrf|| pb_rdf) begin//write_through or read first
        if(cfg_b[3:0]== 4'b1100 || cfg_b[3:0]== 4'b1110 || cfg_b[3:0]== 4'b1111) begin
        do_b={2'bx,do_b_comb[15:0]};
        end
        else begin
        do_b=do_b_comb;
        end
      end	  
      else begin // write no-change mode
       do_b=do_b ;
      end
    end
  end
// else if (~por_b) do_b=0;
end	    
endmodule
//FIFO Controller Core
`ifndef DLY
`define DLY #1
`endif

module fifo_ctrl_core(
		w_width,
		r_width,
		depth_ext_mode,
		peek_mode,
		wclk,
		rclk,
		wrst_n,
		rrst_n,
		wr_req_n,
		write_drop,
		write_save,
		wrdp_rd_flag,
		rd_req_n,
		full,
		empty,
		prog_full,
		usr_pf,
		prog_empty,
		usr_pe,
		overflow,
		underflow,
		wr_mem_n,
		rd_mem_n,
		wr_addr,
		rd_addr
		);

parameter ASIZE		=	14;//address width

input	[3:0]		w_width;
input	[3:0]		r_width;
input	[1:0]		depth_ext_mode;//other for 4.5k, 01 for 9k, 11 for 18k?
input				peek_mode;
input				wclk;
input				rclk;
input				wrst_n;
input				rrst_n;
input				wr_req_n;
input				write_drop;
input				write_save;
input				rd_req_n;
input	[ASIZE-1:0]	usr_pf;//user defined programmable-full level
input	[ASIZE-1:0]	usr_pe;//user defined programmable-empty level

output				full;
output				empty;
output				prog_full;
output				prog_empty;
output				overflow;
output				underflow;
output				wr_mem_n;
output				rd_mem_n;
output	[ASIZE-1:0]	wr_addr;
output	[ASIZE-1:0]	rd_addr;
output				wrdp_rd_flag;

reg					wrdp_rd_flag;
wire				wrdp_rd_jj;
reg					wr_return;
reg					rd_return;
reg					wr_ack;
reg					rd_ack;
reg					overflow;
reg					underflow;

wire	[ASIZE-1:0]	wr_addr;//binary-code address
wire	[ASIZE-1:0]	rd_addr;
wire	[ASIZE-1:0]	wr_gray;//gray-code
wire	[ASIZE-1:0]	rd_gray;
wire	[ASIZE-1:0]	wr_bptr_mask;
wire	[ASIZE-1:0]	rd_bptr_mask;
reg		[ASIZE-1:0]	wr2rd_gray,wr2rd_gray_t;
reg		[ASIZE-1:0]	rd2wr_gray,rd2wr_gray_t;
reg		[ASIZE-1:0]	waddr_save;//for write drop function 
wire	[ASIZE-1:0]	rd2wr_bin;
wire	[ASIZE-1:0]	wr2rd_bin;
reg		[ASIZE-1:0]	wr_bptr;//binary-code
reg		[ASIZE-1:0]	wr_bptr_dly;
reg		[ASIZE-1:0]	rd_bptr;
reg		[ASIZE-1:0]	rd_bptr_dly;
wire				wr_mem_n;
wire				rd_mem_n;
wire	[ASIZE-1:0]	max_step;
wire				wr_rd_diff;//1 : write step gt read step, 0 : read gt write
reg					full;
reg					empty;
reg					full_pre0,full_pre1;
reg					empty_pre0,empty_pre1,empty_pre2;
wire				full_flag;
wire				empty_flag;
wire				wamax;
wire				ramax;
wire	[2:0]		shiftw,shiftr,shift_diff;
wire	[ASIZE:0]	depth,w_depth,r_depth;
wire				gt;

assign depth = 1 << ASIZE;//max fifo depth
//write & read step definition. based on data width.
assign w_depth =	(depth_ext_mode == 2'b11) ? (w_width[0] ? depth					:
												 w_width[1] ? {1'b0,depth[ASIZE:1]} :
												 w_width[2] ? {2'b0,depth[ASIZE:2]} :
												 w_width[3] ? {3'b0,depth[ASIZE:3]} : {4'b0,depth[ASIZE:4]}):
					(depth_ext_mode == 2'b01) ? (w_width[0] ? {1'b0,depth[ASIZE:1]} :
												 w_width[1] ? {2'b0,depth[ASIZE:2]} :
												 w_width[2] ? {3'b0,depth[ASIZE:3]} :
												 w_width[3] ? {4'b0,depth[ASIZE:4]} : {5'b0,depth[ASIZE:5]}):
												(w_width[0] ? {2'b0,depth[ASIZE:2]} :
												 w_width[1] ? {3'b0,depth[ASIZE:3]} :
                                                 w_width[2] ? {4'b0,depth[ASIZE:4]} :
                                                 w_width[3] ? {5'b0,depth[ASIZE:5]} : {6'b0,depth[ASIZE:6]});



assign r_depth = wr_rd_diff ? (w_depth << shift_diff) : (w_depth >> shift_diff);
assign shiftw = w_width[0] ? 0 :
				w_width[1] ? 1 :
				w_width[2] ? 2 :
				w_width[3] ? 3 : 4;
assign shiftr = r_width[0] ? 0 :
				r_width[1] ? 1 :
				r_width[2] ? 2 :
				r_width[3] ? 3 : 4;
assign shift_diff = (shiftw >= shiftr) ? (shiftw - shiftr) : (shiftr - shiftw);
assign max_step = (shiftw >= shiftr) ? shiftw : shiftr;
assign wr_rd_diff = (shiftw >= shiftr) ? 1 : 0;

//write pointer INC & write pointer delay
always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0)	wr_bptr_dly <= `DLY 0;
	else if(write_drop == 1) wr_bptr_dly <= `DLY waddr_save;
	else if(wr_req_n == 0 && full != 1) wr_bptr_dly <= `DLY wr_bptr;
end
always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) wr_bptr <= `DLY 1;
	else if(write_drop == 1) wr_bptr <= `DLY waddr_save + 1;
	else if(wr_req_n == 0 && full != 1) wr_bptr <= `DLY wr_bptr + 1;
end
assign wr_addr = (depth_ext_mode == 2'b11) ? (wr_bptr_dly << shiftw) : (depth_ext_mode == 2'b01) ? {1'b0,(wr_bptr_dly[ASIZE-2:0] << shiftw)} : {2'b00,(wr_bptr_dly[ASIZE-3:0] << shiftw)};

//write drop function realization
always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) waddr_save <= `DLY 14'h3fff;
	else if(write_save == 1) waddr_save <= `DLY wr_bptr_dly;
end

//read pointer INC & read pointer delay
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) rd_bptr_dly <= `DLY 0;
	else if(rd_req_n == 0 && empty != 1) rd_bptr_dly <= `DLY rd_bptr;
end
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) begin rd_bptr <= `DLY 1; end
	else if(rd_req_n == 0 && empty != 1) begin rd_bptr <= `DLY rd_bptr + 1; end
end
assign rd_addr = (depth_ext_mode == 2'b11) ? (rd_bptr_dly << shiftr) : (depth_ext_mode == 2'b01) ? {1'b0,(rd_bptr_dly[ASIZE-2:0] << shiftr)} : {2'b00,(rd_bptr_dly[ASIZE-3:0] << shiftr)};

//binary pointer convert to gray-code
assign wr_bptr_mask =	w_width[0] ? ((depth_ext_mode == 2'b11) ? wr_bptr_dly : (depth_ext_mode == 2'b01) ? {1'b0,wr_bptr_dly[ASIZE-2:0]} : {2'b0,wr_bptr_dly[ASIZE-3:0]}) :
						w_width[1] ? ((depth_ext_mode == 2'b11) ? {1'b0,wr_bptr_dly[ASIZE-2:0]} : (depth_ext_mode == 2'b01) ? {2'b0,wr_bptr_dly[ASIZE-3:0]} : {3'b0,wr_bptr_dly[ASIZE-4:0]}) :
						w_width[2] ? ((depth_ext_mode == 2'b11) ? {2'b0,wr_bptr_dly[ASIZE-3:0]} : (depth_ext_mode == 2'b01) ? {3'b0,wr_bptr_dly[ASIZE-4:0]} : {4'b0,wr_bptr_dly[ASIZE-5:0]}) :
						w_width[3] ? ((depth_ext_mode == 2'b11) ? {3'b0,wr_bptr_dly[ASIZE-4:0]} : (depth_ext_mode == 2'b01) ? {4'b0,wr_bptr_dly[ASIZE-5:0]} : {5'b0,wr_bptr_dly[ASIZE-6:0]}) :
						((depth_ext_mode == 2'b11) ? {4'b0,wr_bptr_dly[ASIZE-5:0]} : (depth_ext_mode == 2'b01) ? {5'b0,wr_bptr_dly[ASIZE-6:0]} : {6'b0,wr_bptr_dly[ASIZE-7:0]});
assign rd_bptr_mask =	r_width[0] ? ((depth_ext_mode == 2'b11) ? rd_bptr_dly : (depth_ext_mode == 2'b01) ? {1'b0,rd_bptr_dly[ASIZE-2:0]} : {2'b0,rd_bptr_dly[ASIZE-3:0]}) :
						r_width[1] ? ((depth_ext_mode == 2'b11) ? {1'b0,rd_bptr_dly[ASIZE-2:0]} : (depth_ext_mode == 2'b01) ? {2'b0,rd_bptr_dly[ASIZE-3:0]} : {3'b0,rd_bptr_dly[ASIZE-4:0]}) :
						r_width[2] ? ((depth_ext_mode == 2'b11) ? {2'b0,rd_bptr_dly[ASIZE-3:0]} : (depth_ext_mode == 2'b01) ? {3'b0,rd_bptr_dly[ASIZE-4:0]} : {4'b0,rd_bptr_dly[ASIZE-5:0]}) :
						r_width[3] ? ((depth_ext_mode == 2'b11) ? {3'b0,rd_bptr_dly[ASIZE-4:0]} : (depth_ext_mode == 2'b01) ? {4'b0,rd_bptr_dly[ASIZE-5:0]} : {5'b0,rd_bptr_dly[ASIZE-6:0]}) :
						((depth_ext_mode == 2'b11) ? {4'b0,rd_bptr_dly[ASIZE-5:0]} : (depth_ext_mode == 2'b01) ? {5'b0,rd_bptr_dly[ASIZE-6:0]} : {6'b0,rd_bptr_dly[ASIZE-7:0]});

assign wr_gray = (wr_bptr_mask >> 1) ^ wr_bptr_mask;
assign rd_gray = (rd_bptr_mask >> 1) ^ rd_bptr_mask;
//assign empty_spt_gray = (empty_spt >> 1) ^ empty_spt;

//programmable full & programmalbe empty
//read address - write clock domain synchronization
always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) begin rd2wr_gray <= `DLY 0; rd2wr_gray_t <= `DLY 0;end
	else begin rd2wr_gray <= `DLY rd2wr_gray_t; rd2wr_gray_t <= `DLY rd_gray;end
end
//write address - read clock domain synchronization
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) begin wr2rd_gray <= `DLY 0; wr2rd_gray_t <= `DLY 0;end
	else begin wr2rd_gray <= `DLY wr2rd_gray_t; wr2rd_gray_t <= `DLY wr_gray;end
end

//for empty & full judgement.
assign wamax =	(shiftw == 0) ? ((depth_ext_mode == 2'b11) ? (wr_addr == 'h3fff) : (depth_ext_mode == 2'b01) ? (wr_addr == 'h1fff) : (wr_addr == 'h0fff)) :
				(shiftw == 1) ? ((depth_ext_mode == 2'b11) ? (wr_addr == 'h3ffe) : (depth_ext_mode == 2'b01) ? (wr_addr == 'h1ffe) : (wr_addr == 'h0ffe)) :
				(shiftw == 2) ? ((depth_ext_mode == 2'b11) ? (wr_addr == 'h3ffc) : (depth_ext_mode == 2'b01) ? (wr_addr == 'h1ffc) : (wr_addr == 'h0ffc)) :
				(shiftw == 3) ? ((depth_ext_mode == 2'b11) ? (wr_addr == 'h3ff8) : (depth_ext_mode == 2'b01) ? (wr_addr == 'h1ff8) : (wr_addr == 'h0ff8)) :
									((depth_ext_mode == 2'b11) ? (wr_addr == 'h3ff0) : (depth_ext_mode == 2'b01) ? (wr_addr == 'h1ff0) : (wr_addr == 'h0ff0));
assign ramax =	(shiftr == 0) ? ((depth_ext_mode == 2'b11) ? (rd_addr == 'h3fff) : (depth_ext_mode == 2'b01) ? (rd_addr == 'h1fff) :(rd_addr == 'h0fff)) :
				(shiftr == 1) ? ((depth_ext_mode == 2'b11) ? (rd_addr == 'h3ffe) : (depth_ext_mode == 2'b01) ? (rd_addr == 'h1ffe) : (rd_addr == 'h0ffe)) :
				(shiftr == 2) ? ((depth_ext_mode == 2'b11) ? (rd_addr == 'h3ffc) : (depth_ext_mode == 2'b01) ? (rd_addr == 'h1ffc) : (rd_addr == 'h0ffc)) :
				(shiftr == 3) ? ((depth_ext_mode == 2'b11) ? (rd_addr == 'h3ff8) : (depth_ext_mode == 2'b01) ? (rd_addr == 'h1ff8) : (rd_addr == 'h0ff8)) :
									((depth_ext_mode == 2'b11) ? (rd_addr == 'h3ff0) : (depth_ext_mode == 2'b01) ? (rd_addr == 'h1ff0) :(rd_addr == 'h0ff0));


always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) wr_return <= `DLY 0;
	else if(wamax == 1 && wr_req_n == 0 && ~full) wr_return <= `DLY ~wr_return;
end
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) rd_return <= `DLY 0;
	else if(ramax == 1 && rd_req_n == 0 && ~empty) rd_return <= `DLY ~rd_return;
end

assign gt = (wr_return == rd_return) ? 1 : 0;

//memory control signals
assign wr_mem_n = wr_req_n | full;
assign rd_mem_n = rd_req_n | empty;//peek_mode ? empty_pre0 : (rd_req_n | empty);

//full & empty signals generation
assign full_flag = (wr_return != rd_return) && (~empty) && (shift_diff == 0 ? wr_gray == rd_gray : (wr_rd_diff == 1 ? (wr_gray == (rd_gray >> shift_diff)) : (rd_gray == (wr_gray >> shift_diff))));
assign empty_flag = (wr_return == rd_return) && (~full) && (shift_diff == 0 ? wr_gray == rd_gray : (wr_rd_diff == 1 ? (wr_gray == (rd_gray >> shift_diff)) : (rd_gray == (wr_gray >> shift_diff))));

always @(posedge wclk or negedge wrst_n or posedge full_flag)begin
	if(wrst_n == 0) {full,full_pre0,full_pre1} <= `DLY 3'b000;
	else if(full_flag == 1) {full,full_pre0,full_pre1} <= `DLY 3'b111;
	else begin full <= `DLY full_pre0;full_pre0 <= `DLY full_pre1;full_pre1 <= `DLY full_flag;end
end

always @(posedge rclk or negedge rrst_n or posedge empty_flag)begin
	if(rrst_n == 0) {empty,empty_pre0,empty_pre1,empty_pre2} <= `DLY 4'b1111;
	else if(empty_flag == 1) {empty,empty_pre0,empty_pre1,empty_pre2} <= `DLY 4'b1111;
	else begin empty <= `DLY peek_mode ? empty_pre1 : empty_pre0;empty_pre0 <= `DLY empty_pre1;empty_pre1 <= `DLY empty_flag; empty_pre2 <= `DLY empty_flag;end
end

//write drop function read address conflict flag
assign wrdp_rd_jj = (shift_diff == 0 ? waddr_save == rd_bptr_dly : (wr_rd_diff == 1 ? waddr_save == (rd_bptr_dly >> shift_diff) : rd_bptr_dly == (waddr_save >> shift_diff)));
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) wrdp_rd_flag <= `DLY 0;
	else if(wrdp_rd_jj) wrdp_rd_flag <= `DLY 1;
	else if(wrdp_rd_flag == 1 && write_save == 1 && !empty) wrdp_rd_flag <= `DLY 0;
end


//wr_ack & rd_ack signals generation
always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) wr_ack <= `DLY 0;
	else wr_ack <= `DLY (~wr_req_n) & (~full);
end
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) rd_ack <= `DLY 0;
	else rd_ack <= `DLY (~rd_req_n) & (~empty);
end

//overflow & underflow signals generation
always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) overflow <= `DLY 0;
	else overflow <= `DLY (~wr_req_n) & full;
end
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) underflow <= `DLY 0;
	else underflow <= `DLY (~rd_req_n) & empty;
end

gry2bin u0(
	.gry(rd2wr_gray),
	.bin(rd2wr_bin)
	);
gry2bin u1(
	.gry(wr2rd_gray),
	.bin(wr2rd_bin)
	);
prog_fe u2(
	.wclk(wclk),
	.rclk(rclk),
	.wrst_n(wrst_n),
	.rrst_n(rrst_n),
	.prog_full(prog_full),
	.prog_empty(prog_empty),
	.usr_pf(usr_pf),
	.usr_pe(usr_pe),
	.shiftw(shiftw),
	.shiftr(shiftr),
	.depth_ext_mode(depth_ext_mode),
	.wr_addr(wr_bptr_mask),
	.rd_addr(rd_bptr_mask),
	.wr2rd_bin(wr2rd_bin),
	.rd2wr_bin(rd2wr_bin),
	.full(full),
	.empty(empty),
	.w_depth(w_depth),
	.r_depth(r_depth),
	.gt(gt),
	.shift_diff(shift_diff),
	.wr_rd_diff(wr_rd_diff)
	);
endmodule

//gray-code to binary-code transfermation function
module gry2bin(gry,bin);
parameter ASIZE = 14; 
input	[ASIZE-1:0]	gry; 
output	[ASIZE-1:0]	bin; 

reg [ASIZE-1:0] bin; 
integer i;
always @(gry)
begin    
    bin[ASIZE-1]=gry[ASIZE-1];    
    for(i=ASIZE-2;i>=0;i=i-1)        
        bin[i]=bin[i+1]^gry[i];
end
endmodule

//programmbale-full & programmable-empty judgement module
module prog_fe(
	wclk,
	rclk,
	wrst_n,
	rrst_n,
	prog_full,
	prog_empty,
	usr_pf,
	usr_pe,
	shiftw,
	shiftr,
	depth_ext_mode,
	wr_addr,
	rd_addr,
	wr2rd_bin,
	rd2wr_bin,
	full,
	empty,
	w_depth,
	r_depth,
	gt,
	shift_diff,
	wr_rd_diff
	);

parameter	ASIZE = 14;
output				prog_full;
output				prog_empty;
input				wclk;//for write full
input				rclk;//for read empty
input				wrst_n;
input				rrst_n;
input	[ASIZE-1:0]	usr_pf;
input	[ASIZE-1:0]	usr_pe;
input	[2:0]		shiftw;
input	[2:0]		shiftr;
input	[1:0]		depth_ext_mode;
input	[ASIZE-1:0]	wr_addr;
input	[ASIZE-1:0]	rd_addr;
input	[ASIZE-1:0]	wr2rd_bin;
input	[ASIZE-1:0]	rd2wr_bin;
input				full;
input				empty;
input	[ASIZE:0]	w_depth;
input	[ASIZE:0]	r_depth;
input				gt;
input	[2:0]		shift_diff;
input				wr_rd_diff;
wire	[ASIZE-1:0]	spt_pf,spt_pe;
wire	[ASIZE-1:0]	rd2wr_s,wr2rd_s;

reg					prog_full;
reg					prog_empty;
wire				cross_pf,cross_pe;

//debug segment//comment out when rtl was frozen

assign rd2wr_s = wr_rd_diff ? (rd2wr_bin >> shift_diff) : (rd2wr_bin << shift_diff);
assign wr2rd_s = wr_rd_diff ? (wr2rd_bin << shift_diff) : (wr2rd_bin >> shift_diff);
assign cross_pf = (rd2wr_s >= wr_addr) ? 0 : 1;
assign cross_pe = (wr2rd_s >= rd_addr) ? 1 : 0;
assign spt_pf = (cross_pf ? w_depth : 0) + rd2wr_s - wr_addr;
assign spt_pe = (cross_pe ? 0 : r_depth) + wr2rd_s - rd_addr;

always @(posedge wclk or negedge wrst_n)begin
	if(wrst_n == 0) prog_full <= `DLY 0;
	else prog_full <= `DLY ((spt_pf <= (usr_pf >> shiftw)) & ~empty) | full;
end
always @(posedge rclk or negedge rrst_n)begin
	if(rrst_n == 0) prog_empty <= `DLY 1;
	else prog_empty <= `DLY ((spt_pe <= (usr_pe >> shiftr)) & ~full) | empty;
end
endmodule
//use in peek-mode to pre-read data from master fifo.
`ifndef DLY
`define DLY #1
`endif

module fifo_pkarbit(
	clk,
	rst_n,
	empty_m,
	full_s,//full & empty from slave fifo
	afull_s,
	rd_n_m,//read require to master fifo
	wr_n_s,//write require to slave fifo
	rd_req_usr //user read require,may be useless too
	);

input			clk;
input			rst_n;
input			empty_m;
input			full_s,afull_s;
input			rd_req_usr;
output			rd_n_m;
output			wr_n_s;

wire			rd_n_m,rd_n_s;
wire			act;
reg				rw_act;
reg				wr_n_s;

assign act = (/*afull_s | */full_s) & rd_req_usr | empty_m;
//assign act = (/*afull_s |*/ full_s | empty_m ) & rd_req_usr;

assign rd_n_m = act;
always @(posedge clk or negedge rst_n)begin
	if(rst_n == 0) wr_n_s <= `DLY 1;
	else wr_n_s <= `DLY act;
end


endmodule


//small module for peek mode.
`ifndef DLY
`define DLY #1
`endif

module fifo_pkslice(
	clk,//write & read use common clock
	rst_n,//common reset
	wr_req_n,
	rd_req_n,
	full,
	afull,
	empty,
	overflow,
	underflow,
	wr_en,
	rd_en
	);

input				clk;
input				rst_n;
input				wr_req_n;
input				rd_req_n;
output				full;
output				afull;
output				empty;
output				overflow;
output				underflow;
output				wr_en;
output				rd_en;

reg					empty,full_i,afull;
reg					overflow,underflow;
reg					wrp,rdp;
wire				full;

always @(posedge clk or negedge rst_n)begin
	if(rst_n == 0) begin
		wrp <= `DLY 0; rdp <= `DLY 0; empty <= `DLY 1; full_i <= `DLY 0; afull <= `DLY 0;
		overflow <= `DLY 0; underflow <= `DLY 0;
		end
	else
		case({wr_req_n,rd_req_n})
			2'b00://write & read at same time
				begin
					if(empty == 1)begin underflow <= `DLY 1; wrp <= `DLY wrp + 1;empty <= `DLY 0;afull <= `DLY 1;end
					else if(full_i == 1)begin overflow <= `DLY 1; rdp <= `DLY rdp + 1;full_i <= `DLY 0;afull <= `DLY 1;underflow <= `DLY 0;end
					else begin wrp <= `DLY wrp + 1; rdp <= `DLY rdp + 1; afull <= `DLY 1;
								underflow <= `DLY 0; overflow <= `DLY 0;end
				end
			2'b01://write only
				begin
					if(full_i == 1)begin overflow <= `DLY 1;end
					else if(wrp != rdp) begin wrp <= `DLY wrp + 1; full_i <= `DLY 1; afull <= `DLY 0; 
												overflow <= `DLY 0;end
					else begin wrp <= `DLY wrp + 1; empty <= `DLY 0; afull <= `DLY 1; overflow <= `DLY 0;end
					underflow <= `DLY 0;
				end
			2'b10://read only
				begin
					if(empty == 1)begin underflow <= `DLY 1;end
					else if(wrp != rdp) begin rdp <= `DLY rdp + 1; empty <= `DLY 1; afull <= `DLY 0; underflow <= `DLY 0;end
					else begin rdp <= `DLY rdp + 1; full_i <= `DLY 0; underflow <= `DLY 0;afull <= 1;end
				end
			2'b11:
				begin
					underflow <= `DLY 0;
					overflow <= `DLY 0;
				end
				//11: no op. and default is a latch
		endcase
end
assign full = full_i | (afull & ~wr_req_n);

assign wr_en = (full_i & rd_req_n) ? ~wrp : wrp;
assign rd_en = empty ? ~rdp : rdp;



endmodule

module glbsr( GSR );

parameter T_GLBSR = 1;

output GSR;
reg GSR_t;

assign (weak1, weak0) GSR = GSR_t;

initial begin
    GSR_t = 1'b0;
    #(T_GLBSR)
    GSR_t = 1'b1;
end

endmodule


module CLK (
	fclk0_il,
	fclk0_oen,
	fclk0_ol,
	fclk1_il,
	fclk1_ol,
	geclk0_il,
	geclk0_ol,
	geclk0_up_il,
	geclk0_up_ol,
	geclk1_il,
	geclk1_ol,
	gsclk0_il,
	gsclk0_ol,
	gsclk1_il,
	gsclk1_ol,
	id_rst,
	id_setn,
	od_rst,
	od_setn,
	oen_rst,
	oen_setn,
	//PARAMETER 
	CFG_CKEN_INV,
	CFG_CKEN_INV_,
	CFG_FCLK0_I_EN,
	CFG_FCLK0_OEN,
	CFG_FCLK0_O_EN,
	CFG_FCLK0_RS_EN,
	CFG_FCLK0_UPI_EN,
	CFG_FCLK0_UPO_EN,
	CFG_FCLK1_I_EN,
	CFG_FCLK1_O_EN,
	CFG_GECLK0_I_EN,
	CFG_GECLK0_O_EN,
	CFG_GECLK1_I_EN,
	CFG_GECLK1_O_EN,
	CFG_GSCLK0_I_EN,
	CFG_GSCLK0_O_EN,
	CFG_GSCLK1_I_EN,
	CFG_GSCLK1_O_EN,
	CFG_RSTN_ID_EN,
	CFG_RSTN_ID_EN_,
	CFG_RSTN_INV,
	CFG_RSTN_INV_,
	CFG_RSTN_OD_EN,
	CFG_RSTN_OD_EN_,
	CFG_RSTN_OEN_EN,
	CFG_RSTN_OEN_EN_,
	CFG_RSTN_SYNC,
	CFG_RSTN_SYNC_,
	CFG_SETN_ID_EN,
	CFG_SETN_ID_EN_,
	CFG_SETN_INV,
	CFG_SETN_INV_,
	CFG_SETN_OD_EN,
	CFG_SETN_OD_EN_,
	CFG_SETN_OEN_EN,
	CFG_SETN_OEN_EN_,
	CFG_SETN_SYNC,
	CFG_SETN_SYNC_,
	CFG_SCLK_INV,
	CFG_ECLK_INV,
	//PARAMETER END
	setn,
	rstn,
	clk_en,
	sclk,
	feclk
	);
output	fclk0_il;
output	fclk0_oen;
output	fclk0_ol;
output	fclk1_il;
output	fclk1_ol;
output	geclk0_il;
output	geclk0_ol;
output	geclk0_up_il;
output	geclk0_up_ol;
output	geclk1_il;
output	geclk1_ol;
output	gsclk0_il;
output	gsclk0_ol;
output	gsclk1_il;
output	gsclk1_ol;
output	id_rst;
output	id_setn;
output	od_rst;
output	od_setn;
output	oen_rst;
output	oen_setn;
input	CFG_CKEN_INV;
input	CFG_CKEN_INV_;
input	CFG_FCLK0_I_EN;
input	CFG_FCLK0_OEN;
input	CFG_FCLK0_O_EN;
input	CFG_FCLK0_RS_EN;
input	CFG_FCLK0_UPI_EN;
input	CFG_FCLK0_UPO_EN;
input	CFG_FCLK1_I_EN;
input	CFG_FCLK1_O_EN;
input	CFG_GECLK0_I_EN;
input	CFG_GECLK0_O_EN;
input	CFG_GECLK1_I_EN;
input	CFG_GECLK1_O_EN;
input	CFG_GSCLK0_I_EN;
input	CFG_GSCLK0_O_EN;
input	CFG_GSCLK1_I_EN;
input	CFG_GSCLK1_O_EN;
input	CFG_RSTN_ID_EN;
input	CFG_RSTN_ID_EN_;
input	CFG_RSTN_INV;
input	CFG_RSTN_INV_;
input	CFG_RSTN_OD_EN;
input	CFG_RSTN_OD_EN_;
input	CFG_RSTN_OEN_EN;
input	CFG_RSTN_OEN_EN_;
input	CFG_RSTN_SYNC;
input	CFG_RSTN_SYNC_;
input	CFG_SETN_ID_EN;
input	CFG_SETN_ID_EN_;
input	CFG_SETN_INV;
input	CFG_SETN_INV_;
input	CFG_SETN_OD_EN;
input	CFG_SETN_OD_EN_;
input	CFG_SETN_OEN_EN;
input	CFG_SETN_OEN_EN_;
input	CFG_SETN_SYNC;
input	CFG_SETN_SYNC_;
input	CFG_SCLK_INV;
input	CFG_ECLK_INV;
input	setn;
input	rstn;
input	clk_en;
input	sclk;
input	feclk;

wire ck_inv = ({CFG_CKEN_INV,CFG_CKEN_INV_} == 2'b01) ? clk_en :
			  ({CFG_CKEN_INV,CFG_CKEN_INV_} == 2'b10) ? ~clk_en : 1'b0;
wire sckinv = CFG_SCLK_INV ? ~sclk  : sclk;
wire eckinv = CFG_ECLK_INV ? ~feclk : feclk;
wire sclk_b,eclk_b;
reg	sck_reg,eck_reg;
always @(sckinv or ck_inv)
	if(sckinv == 0) sck_reg <= ck_inv;
always @(eckinv or ck_inv)
	if(eckinv == 0) eck_reg <= ck_inv;
assign sclk_b = (sckinv & sck_reg);
assign eclk_b = (eckinv & eck_reg);

wire fclk0_sr;
assign fclk0_sr = CFG_FCLK0_RS_EN & eclk_b;
assign geclk0_up_il = CFG_FCLK0_UPI_EN & eclk_b;
assign geclk0_up_ol = CFG_FCLK0_UPO_EN & eclk_b;
assign fclk0_oen = CFG_FCLK0_OEN & eclk_b;
assign geclk0_il = CFG_GECLK0_I_EN & eclk_b;
assign geclk1_il = CFG_GECLK1_I_EN & eclk_b;
assign fclk0_il = CFG_FCLK0_I_EN & eclk_b;
assign fclk1_il = CFG_FCLK1_I_EN & eclk_b;
assign geclk0_ol = CFG_GECLK0_O_EN & eclk_b;
assign geclk1_ol = CFG_GECLK1_O_EN & eclk_b;
assign fclk0_ol = CFG_FCLK0_O_EN & eclk_b;
assign fclk1_ol = CFG_FCLK1_O_EN & eclk_b;
assign gsclk0_ol = CFG_GSCLK0_O_EN & sclk_b;
assign gsclk1_ol = CFG_GSCLK1_O_EN & sclk_b;
assign gsclk0_il = CFG_GSCLK0_I_EN & sclk_b;
assign gsclk1_il = CFG_GSCLK1_I_EN & sclk_b;

wire set_inv = ({CFG_SETN_INV,CFG_SETN_INV_} == 2'b01) ? ~setn :
			   ({CFG_SETN_INV,CFG_SETN_INV_} == 2'b10) ? setn : 1'b0;
reg	set_reg;
always @(set_inv or fclk0_sr)
	if(fclk0_sr == 0) set_reg <= set_inv;
wire set_sync = (set_reg & fclk0_sr);
wire set_sel = ({CFG_SETN_SYNC,CFG_SETN_SYNC_} == 2'b01) ? set_inv :
			   ({CFG_SETN_SYNC,CFG_SETN_SYNC_} == 2'b10) ? set_sync : 1'b0;
wire od_set = ({CFG_SETN_OD_EN,CFG_SETN_OD_EN_} == 2'b01) ? 1'b1 :
			  ({CFG_SETN_OD_EN,CFG_SETN_OD_EN_} == 2'b10) ? ~set_sel : 1'b0;
wire id_set = ({CFG_SETN_ID_EN,CFG_SETN_ID_EN_} == 2'b01) ? 1'b1 :
			  ({CFG_SETN_ID_EN,CFG_SETN_ID_EN_} == 2'b10) ? ~set_sel : 1'b0;
wire oen_set = ({CFG_SETN_OEN_EN,CFG_SETN_OEN_EN_} == 2'b01) ? 1'b1 :
			   ({CFG_SETN_OEN_EN,CFG_SETN_OEN_EN_} == 2'b10) ? ~set_sel : 1'b0;
assign od_setn = od_set;
assign id_setn = id_set;
assign oen_setn = oen_set;
wire rst_inv = ({CFG_RSTN_INV,CFG_RSTN_INV_} == 2'b01) ? ~rstn :
			   ({CFG_RSTN_INV,CFG_RSTN_INV_} == 2'b10) ? rstn : 1'b0;
reg	rst_reg;
always @(rst_inv or fclk0_sr)
	if(fclk0_sr == 0) rst_reg <= rst_inv;
wire rst_sync = (rst_reg & fclk0_sr);
wire rst_sel = ({CFG_RSTN_SYNC,CFG_RSTN_SYNC_} == 2'b01) ? rst_inv :
			   ({CFG_RSTN_SYNC,CFG_RSTN_SYNC_} == 2'b10) ? rst_sync : 1'b0;
wire od_rst = ({CFG_RSTN_OD_EN,CFG_RSTN_OD_EN_} == 2'b01) ? 1'b0 :
			  ({CFG_RSTN_OD_EN,CFG_RSTN_OD_EN_} == 2'b10) ? rst_sel : 1'b1;
wire id_rst = ({CFG_RSTN_ID_EN,CFG_RSTN_ID_EN_} == 2'b01) ? 1'b0 :
			  ({CFG_RSTN_ID_EN,CFG_RSTN_ID_EN_} == 2'b10) ? rst_sel : 1'b1;
wire oen_rst = ({CFG_RSTN_OEN_EN,CFG_RSTN_OEN_EN_} == 2'b01) ? 1'b0 :
			   ({CFG_RSTN_OEN_EN,CFG_RSTN_OEN_EN_} == 2'b10) ? rst_sel : 1'b1;

endmodule

module ILOGIC (
	//in & out
	shiftout0,
	shiftout1,
	dataout,

	datain,
	fclk0,
	fclk1,
	geclk0,
	geclk1,
	gsclk0,
	gsclk1,
	init_b,
	rst,
	set_,
	shiftin0,
	shiftin1,
	update,
	update_,
	usermode,
	test,
	//parameter
	CFG_DDR_IN_NREG,
	CFG_DDR_IN_NREG_DFF,
	CFG_DDR_IN_PREG,
	CFG_DDR_IN_PREG_DFF,
	CFG_DQS_CLK,
	CFG_FASTIN,
	CFG_SLAVE_IN,
	CFG_TEST,
	CFG_IN_EN,
	CFG_GEAR_IN,
	CFG_DDR_IN_NREG_,
	CFG_DDR_IN_NREG_DFF_,
	CFG_DDR_IN_PREG_,
	CFG_DDR_IN_PREG_DFF_,
	CFG_DQS_CLK_,
	CFG_FASTIN_,
	CFG_SLAVE_IN_,
	CFG_TEST_,
	CFG_IN_EN_,
	CFG_GEAR_IN_
	);
output	shiftout0,shiftout1;
output	[7:0]	dataout;
input	datain;
input	fclk0;
input	fclk1;
input	geclk0;
input	geclk1;
input	gsclk0;
input	gsclk1;
input	init_b;
input	rst;
input	set_;
input	shiftin0;
input	shiftin1;
input	update,update_;
input	usermode;
input	[7:0]	test;

input	CFG_DDR_IN_NREG;
input	CFG_DDR_IN_NREG_DFF;
input	CFG_DDR_IN_PREG;
input	CFG_DDR_IN_PREG_DFF;
input	CFG_DQS_CLK;
input	CFG_FASTIN;
input	CFG_SLAVE_IN;
input	[7:0]	CFG_TEST;
input	[1:0]	CFG_IN_EN;
input	[7:0]	CFG_GEAR_IN;
input	CFG_DDR_IN_NREG_;
input	CFG_DDR_IN_NREG_DFF_;
input	CFG_DDR_IN_PREG_;
input	CFG_DDR_IN_PREG_DFF_;
input	CFG_DQS_CLK_;
input	CFG_FASTIN_;
input	CFG_SLAVE_IN_;
input	[7:0]	CFG_TEST_;
input	[1:0]	CFG_IN_EN_;
input	[7:0]	CFG_GEAR_IN_;

wire	usermode_b=~usermode;
wire	clk_n,clk_p;
assign clk_n = ({CFG_DQS_CLK,CFG_DQS_CLK_} == 2'b01) ? fclk1 :
			   ({CFG_DQS_CLK,CFG_DQS_CLK_} == 2'b10) ? 1'b1 : 1'bx;
assign clk_p = ({CFG_DQS_CLK,CFG_DQS_CLK_} == 2'b01) ? ~fclk0 :
			   ({CFG_DQS_CLK,CFG_DQS_CLK_} == 2'b10) ? 1'b1 : 1'bx;
reg		nreg_n,nreg_p;//clk_n path register. active @ negedge/posedge
reg		preg_n,preg_n2;//clk_p path register are all active @ negedge of clk_p
always @(negedge clk_n or posedge rst or negedge set_)
	if(set_ == 0) nreg_n <= 1;
	else if(rst) nreg_n <= 0;
	else nreg_n <= datain;
always @(posedge clk_n or posedge rst or negedge set_)
	if(set_ == 0) nreg_p <= 1;
	else if(rst) nreg_p <= 0;
	else nreg_p <= nreg_n;
always @(negedge clk_p or posedge rst or negedge set_)
	if(set_ == 0) preg_n <= 1;
	else if(rst) preg_n <= 0;
	else preg_n <= datain;
always @(negedge clk_p or posedge rst or negedge set_)
	if(set_ == 0) preg_n2 <= 1;
	else if(rst) preg_n2 <= 0;
	else preg_n2 <= preg_n;

wire	n_sel,p_sel;
assign n_sel =	({CFG_FASTIN,CFG_DDR_IN_NREG,CFG_DDR_IN_NREG_DFF,CFG_FASTIN_,CFG_DDR_IN_NREG_,CFG_DDR_IN_NREG_DFF_} == 6'b100011) ? datain :
				({CFG_FASTIN,CFG_DDR_IN_NREG,CFG_DDR_IN_NREG_DFF,CFG_FASTIN_,CFG_DDR_IN_NREG_,CFG_DDR_IN_NREG_DFF_} == 6'b010101) ? nreg_n :
				({CFG_FASTIN,CFG_DDR_IN_NREG,CFG_DDR_IN_NREG_DFF,CFG_FASTIN_,CFG_DDR_IN_NREG_,CFG_DDR_IN_NREG_DFF_} == 6'b001110) ? nreg_p :
				({CFG_FASTIN,CFG_DDR_IN_NREG,CFG_DDR_IN_NREG_DFF,CFG_FASTIN_,CFG_DDR_IN_NREG_,CFG_DDR_IN_NREG_DFF_} == 6'b000111) ? 1'b1 : 1'bx;
assign p_sel =	({CFG_FASTIN,CFG_DDR_IN_PREG,CFG_DDR_IN_PREG_DFF,CFG_FASTIN_,CFG_DDR_IN_PREG_,CFG_DDR_IN_PREG_DFF_} == 6'b100011) ? datain :
				({CFG_FASTIN,CFG_DDR_IN_PREG,CFG_DDR_IN_PREG_DFF,CFG_FASTIN_,CFG_DDR_IN_PREG_,CFG_DDR_IN_PREG_DFF_} == 6'b010101) ? preg_n :
				({CFG_FASTIN,CFG_DDR_IN_PREG,CFG_DDR_IN_PREG_DFF,CFG_FASTIN_,CFG_DDR_IN_PREG_,CFG_DDR_IN_PREG_DFF_} == 6'b001110) ? preg_n2 :
				({CFG_FASTIN,CFG_DDR_IN_PREG,CFG_DDR_IN_PREG_DFF,CFG_FASTIN_,CFG_DDR_IN_PREG_,CFG_DDR_IN_PREG_DFF_} == 6'b000111) ? 1'b1 : 1'bx;
reg	q5,q3,q1;//geclk1,clk_n
reg	q4,q2,q0;//geclk0,clk_p
wire	q7,q6;
dff_n2mx q7mx(.q(q7),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(CFG_SLAVE_IN),.sel_(CFG_SLAVE_IN_),.init_b(init_b),.in0(n_sel),.in1(shiftin1));
dff_n2mx q6mx(.q(q6),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(CFG_SLAVE_IN),.sel_(CFG_SLAVE_IN_),.init_b(init_b),.in0(p_sel),.in1(shiftin0));
always @(posedge geclk1 or negedge usermode)begin
	if(~usermode) q5 <= 1;
	else q5 <= q7;
end
always @(posedge geclk0 or negedge usermode)begin
	if(~usermode) q4 <= 1;
	else q4 <= q6;
end
always @(posedge geclk1 or negedge usermode)begin
	if(~usermode) q3 <= 1;
	else q3 <= q5;
end
always @(posedge geclk0 or negedge usermode)begin
	if(~usermode) q2 <= 1;
	else q2 <= q4;
end
always @(posedge geclk1 or negedge usermode)begin
	if(~usermode) q1 <= 1;
	else q1 <= q3;
end
always @(posedge geclk0 or negedge usermode)begin
	if(~usermode) q0 <= 1;
	else q0 <= q2;
end

wire q7s,q5s,q3s,q1s;//update register. active by geclk1
wire q6s,q4s,q2s,q0s;//update register. active by geclk0
dff_2mx q7smx(.q(q7s),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q7s),.in1(q7));
dff_2mx q6smx(.q(q6s),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q6s),.in1(q6));
dff_2mx q5smx(.q(q5s),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q5s),.in1(q5));
dff_2mx q4smx(.q(q4s),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q4s),.in1(q4));
dff_2mx q3smx(.q(q3s),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q3s),.in1(q3));
dff_2mx q2smx(.q(q2s),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q2s),.in1(q2));
dff_2mx q1smx(.q(q1s),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q1s),.in1(q1));
dff_2mx q0smx(.q(q0s),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(q0s),.in1(q0));

reg q7e,q5e,q3e,q1e;//gsclk sync register. active by gsclk1
reg q6e,q4e,q2e,q0e;//gsclk sync register. active by gsclk0
always @(posedge gsclk1 or negedge usermode)begin
	if(~usermode) q7e <= 1;
	else q7e <= q7s;
end
always @(posedge gsclk0 or negedge usermode)begin
	if(~usermode) q6e <= 1;
	else q6e <= q6s;
end
always @(posedge gsclk1 or negedge usermode)begin
	if(~usermode) q5e <= 1;
	else q5e <= q5s;
end
always @(posedge gsclk0 or negedge usermode)begin
	if(~usermode) q4e <= 1;
	else q4e <= q4s;
end
always @(posedge gsclk1 or negedge usermode)begin
	if(~usermode) q3e <= 1;
	else q3e <= q3s;
end
always @(posedge gsclk0 or negedge usermode)begin
	if(~usermode) q2e <= 1;
	else q2e <= q2s;
end
always @(posedge gsclk1 or negedge usermode)begin
	if(~usermode) q1e <= 1;
	else q1e <= q1s;
end
always @(posedge gsclk0 or negedge usermode)begin
	if(~usermode) q0e <= 1;
	else q0e <= q0s;
end

assign dataout[7] =	({CFG_GEAR_IN[7],CFG_TEST[7],CFG_GEAR_IN_[7],CFG_TEST_[7]} == 4'b0110) ? test[7] :
					({CFG_GEAR_IN[7],CFG_TEST[7],CFG_GEAR_IN_[7],CFG_TEST_[7]} == 4'b1001) ? q7e :
					({CFG_GEAR_IN[7],CFG_TEST[7],CFG_GEAR_IN_[7],CFG_TEST_[7]} == 4'b0011) ? 1'b1 : 1'bx;
assign dataout[6] =	({CFG_GEAR_IN[6],CFG_TEST[6],CFG_GEAR_IN_[6],CFG_TEST_[6]} == 4'b0110) ? test[6] :
					({CFG_GEAR_IN[6],CFG_TEST[6],CFG_GEAR_IN_[6],CFG_TEST_[6]} == 4'b1001) ? q6e :
					({CFG_GEAR_IN[6],CFG_TEST[6],CFG_GEAR_IN_[6],CFG_TEST_[6]} == 4'b0011) ? 1'b1 : 1'bx;
assign dataout[5] =	({CFG_GEAR_IN[5],CFG_TEST[5],CFG_GEAR_IN_[5],CFG_TEST_[5]} == 4'b0110) ? test[5] :
					({CFG_GEAR_IN[5],CFG_TEST[5],CFG_GEAR_IN_[5],CFG_TEST_[5]} == 4'b1001) ? q5e :
					({CFG_GEAR_IN[5],CFG_TEST[5],CFG_GEAR_IN_[5],CFG_TEST_[5]} == 4'b0011) ? 1'b1 : 1'bx;
assign dataout[4] =	({CFG_GEAR_IN[4],CFG_TEST[4],CFG_GEAR_IN_[4],CFG_TEST_[4]} == 4'b0110) ? test[4] :
					({CFG_GEAR_IN[4],CFG_TEST[4],CFG_GEAR_IN_[4],CFG_TEST_[4]} == 4'b1001) ? q4e :
					({CFG_GEAR_IN[4],CFG_TEST[4],CFG_GEAR_IN_[4],CFG_TEST_[4]} == 4'b0011) ? 1'b1 : 1'bx;
assign dataout[3] =	({CFG_GEAR_IN[3],CFG_TEST[3],CFG_GEAR_IN_[3],CFG_TEST_[3]} == 4'b0110) ? test[3] :
					({CFG_GEAR_IN[3],CFG_TEST[3],CFG_GEAR_IN_[3],CFG_TEST_[3]} == 4'b1001) ? q3e :
					({CFG_GEAR_IN[3],CFG_TEST[3],CFG_GEAR_IN_[3],CFG_TEST_[3]} == 4'b0011) ? 1'b1 : 1'bx;
assign dataout[2] =	({CFG_GEAR_IN[2],CFG_TEST[2],CFG_GEAR_IN_[2],CFG_TEST_[2]} == 4'b0110) ? test[2] :
					({CFG_GEAR_IN[2],CFG_TEST[2],CFG_GEAR_IN_[2],CFG_TEST_[2]} == 4'b1001) ? q2e :
					({CFG_GEAR_IN[2],CFG_TEST[2],CFG_GEAR_IN_[2],CFG_TEST_[2]} == 4'b0011) ? 1'b1 : 1'bx;
assign dataout[1] =	({CFG_IN_EN[1],CFG_GEAR_IN[1],CFG_TEST[1],CFG_IN_EN_[1],CFG_GEAR_IN_[1],CFG_TEST_[1]} == 6'b100011) ? n_sel :
					({CFG_IN_EN[1],CFG_GEAR_IN[1],CFG_TEST[1],CFG_IN_EN_[1],CFG_GEAR_IN_[1],CFG_TEST_[1]} == 6'b010101) ? q1e :
					({CFG_IN_EN[1],CFG_GEAR_IN[1],CFG_TEST[1],CFG_IN_EN_[1],CFG_GEAR_IN_[1],CFG_TEST_[1]} == 6'b001110) ? test[1] :
					({CFG_IN_EN[1],CFG_GEAR_IN[1],CFG_TEST[1],CFG_IN_EN_[1],CFG_GEAR_IN_[1],CFG_TEST_[1]} == 6'b000111) ? 1'b1 : 1'bx;
assign dataout[0] =	({CFG_IN_EN[0],CFG_GEAR_IN[0],CFG_TEST[0],CFG_IN_EN_[0],CFG_GEAR_IN_[0],CFG_TEST_[0]} == 6'b100011) ? p_sel :
					({CFG_IN_EN[0],CFG_GEAR_IN[0],CFG_TEST[0],CFG_IN_EN_[0],CFG_GEAR_IN_[0],CFG_TEST_[0]} == 6'b010101) ? q0e :
					({CFG_IN_EN[0],CFG_GEAR_IN[0],CFG_TEST[0],CFG_IN_EN_[0],CFG_GEAR_IN_[0],CFG_TEST_[0]} == 6'b001110) ? test[0] :
					({CFG_IN_EN[0],CFG_GEAR_IN[0],CFG_TEST[0],CFG_IN_EN_[0],CFG_GEAR_IN_[0],CFG_TEST_[0]} == 6'b000111) ? 1'b1 : 1'bx;
assign shiftout1 = q1;
assign shiftout0 = q0;

endmodule

module OLOGIC (
	//data port
	dataout,
	shiftout0,
	shiftout1,

	fclk0,
	fclk1,
	geclk0,
	geclk1,
	gsclk0,
	gsclk1,
	rst,
	set_,
	shiftin0,
	shiftin1,
	update,
	update_,
	usermode,
	datain,
	//PARAMETER
	CFG_DDR_OUT,
	CFG_DDR_OUT_REG,
	CFG_DDR_OUT_REG_,
	CFG_FCLK_INV,
	CFG_FOUT_SEL,
	CFG_FOUT_SEL_,
	CFG_GEAR_OUT,
	CFG_GEAR_OUT_
	);
output	dataout;
output	shiftout0;
output	shiftout1;

input	fclk0;
input	fclk1;
input	geclk0;
input	geclk1;
input	gsclk0;
input	gsclk1;
input	rst;
input	set_;
input	shiftin0;
input	shiftin1;
input	update;
input	update_;
input	usermode;
input	[7:0]	datain;
input	CFG_DDR_OUT;
input	CFG_DDR_OUT_REG;
input	CFG_DDR_OUT_REG_;
input	CFG_FCLK_INV;
input	CFG_FOUT_SEL;
input	CFG_FOUT_SEL_;
input	CFG_GEAR_OUT;
input	CFG_GEAR_OUT_;

wire	usermode_b = ~usermode;
reg	q6,q4,q2,q0;//gsclk0 drive data reg
reg	q7,q5,q3,q1;//gsclk1 drive data reg
wire	s6,s4,s2,s0;//geclk0 drive mux-2 out
wire	s7,s5,s3,s1;//geclk1 drive mux-2 out

always @(posedge gsclk0 or negedge usermode)
	if(~usermode) q6 <= 1;
	else q6 <= datain[6];
always @(posedge gsclk1 or negedge usermode)
	if(~usermode) q7 <= 1;
	else q7 <= datain[7];
always @(posedge gsclk0 or negedge usermode)
	if(~usermode) q4 <= 1;
	else q4 <= datain[4];
always @(posedge gsclk1 or negedge usermode)
	if(~usermode) q5 <= 1;
	else q5 <= datain[5];
always @(posedge gsclk0 or negedge usermode)
	if(~usermode) q2 <= 1;
	else q2 <= datain[2];
always @(posedge gsclk1 or negedge usermode)
	if(~usermode) q3 <= 1;
	else q3 <= datain[3];
always @(posedge gsclk0 or negedge usermode)
	if(~usermode) q0 <= 1;
	else q0 <= datain[0];
always @(posedge gsclk1 or negedge usermode)
	if(~usermode) q1 <= 1;
	else q1 <= datain[1];

dff_2mx s6mx(.q(s6),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(shiftin0),.in1(q6));
dff_2mx s7mx(.q(s7),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(shiftin1),.in1(q7));
dff_2mx s4mx(.q(s4),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(s6),.in1(q4));
dff_2mx s5mx(.q(s5),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(s7),.in1(q5));
dff_2mx s2mx(.q(s2),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(s4),.in1(q2));
dff_2mx s3mx(.q(s3),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(s5),.in1(q3));
dff_2mx s0mx(.q(s0),.clk(geclk0),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(s2),.in1(q0));
dff_2mx s1mx(.q(s1),.clk(geclk1),.set_(1'b1),.rst(usermode_b),.sel(update),.sel_(update_),.in0(s3),.in1(q1));

assign shiftout0 = s0;
assign shiftout1 = s1;

wire	dp_0,dn_0,dp_2,dn_2;
assign dp_0 =	({CFG_GEAR_OUT,CFG_GEAR_OUT_} == 2'b01) ? ~datain[0] :
				({CFG_GEAR_OUT,CFG_GEAR_OUT_} == 2'b10) ? ~s0 : 1'bx;
assign dn_0 =	({CFG_GEAR_OUT,CFG_GEAR_OUT_} == 2'b01) ? ~datain[1] :
				({CFG_GEAR_OUT,CFG_GEAR_OUT_} == 2'b10) ? ~s1 : 1'bx;
reg	dp_1,dp_3;//fclk0 drive
reg	dn_1,dn_3;//fclk1 drive

always @(posedge fclk0 or posedge rst or negedge set_)
	if(~set_) dp_1 <= 1;
	else if(rst) dp_1 <= 0;
	else dp_1 <= dp_0;
always @(posedge fclk1 or posedge rst or negedge set_)
	if(~set_) dn_1 <= 1;
	else if(rst) dn_1 <= 0;
	else dn_1 <= dn_0;

assign dp_2 =	({CFG_DDR_OUT_REG,CFG_DDR_OUT_REG_} == 2'b01) ? ~dp_0 :
				({CFG_DDR_OUT_REG,CFG_DDR_OUT_REG_} == 2'b10) ? ~dp_1 : 1'bx;
assign dn_2 =	({CFG_DDR_OUT_REG,CFG_DDR_OUT_REG_} == 2'b01) ? ~dn_0 :
				({CFG_DDR_OUT_REG,CFG_DDR_OUT_REG_} == 2'b10) ? ~dn_1 : 1'bx;

always @(posedge fclk0 or posedge rst or negedge set_)
	if(~set_) dp_3 <= 1;
	else if(rst) dp_3 <= 0;
	else dp_3 <= dp_2;
always @(negedge fclk1 or posedge rst or negedge set_)
	if(~set_) dn_3 <= 1;
	else if(rst) dn_3 <= 0;
	else dn_3 <= dn_2;

wire	fclk_ddr;
assign fclk_ddr = !(fclk0 & CFG_DDR_OUT);
wire	ck_s_d,ck_s_d_b;
assign ck_s_d = fclk_ddr & CFG_FCLK_INV;
assign ck_s_d_b = !(fclk_ddr & CFG_FCLK_INV);

wire	dp_out;
assign dp_out =	({ck_s_d,ck_s_d_b} == 2'b01) ? dn_3:
				({ck_s_d,ck_s_d_b} == 2'b10) ? dp_3:1'bx;
assign dataout =	({CFG_FOUT_SEL,CFG_FOUT_SEL_} == 2'b01) ? dp_out:
					({CFG_FOUT_SEL,CFG_FOUT_SEL_} == 2'b10) ? datain[0]:1'bx;



endmodule


`ifndef DLY
    `define DLY #1
`endif

module ioc_latn_ar(
     ck
    ,d
    ,q
    ,rstn
);

input  ck;
input  d;
output q;
input  rstn;

reg q;

always@(*)
begin
    if(~rstn)
        q <= `DLY 1'b0;
    else if(ck == 1'b0)
        q <= `DLY d;
end

endmodule

module ioc_dff_asr(
     ck
    ,d
    ,q
    ,rstn
    ,setn
);

input  ck;
input  d;
output q;
input  rstn;
input  setn;

reg q;

always@(posedge ck or negedge setn or negedge rstn)
begin
    if(~rstn)
	q <= `DLY 1'b0;
    else if(~setn)
	q <= `DLY 1'b1;
    else
	q <= `DLY d;
end

endmodule

module ioc_dffn_asr(
     ckb
    ,d
    ,q
    ,rstn
    ,setn
);

input  ckb;
input  d;
output q;
input  rstn;
input  setn;

reg q;

always@(negedge ckb or negedge setn or negedge rstn)
begin
    if(~rstn)
	q <= `DLY 1'b0;
    else if(~setn)
	q <= `DLY 1'b1;
    else
	q <= `DLY d;
end

endmodule


`ifndef CS_SW_SKEL
//----------------------------------------------------------------------------
//
// module: LUT5
//
// description: 5 input lookup-table
// config:      32 bit init value
//
//----------------------------------------------------------------------------
module LUT5 (
         dx,
         f4,
         f3,
         f2,
         f1,
         f0
`ifdef FM_HACK
        ,config_data
`endif
         );

    input       f4;
    input       f3;
    input       f2;
    input       f1;
    input       f0;

    output      dx;

`ifdef CS_FORMALPRO_HACK
    wire [31:0]         config_data;
`else
     `ifdef  SIMULATION
          reg [31:0] config_data = 32'h00000000;
     `else
        `ifdef FM_HACK
            input   [31:0]  config_data;
        `else
            parameter  config_data = 32'h00000000;
        `endif
     `endif
`endif

`ifndef CS_SW_SKEL
    wire [31:0]         cfg = config_data;
    wire [15:0]         da;
    wire [7:0]          db;
    wire [3:0]          dc;
    wire [1:0]          dd;
    wire                de;

    MUX2S_L muxa0(.o(da[0]),  .sel(f0), .i1(cfg[1]), .i0(cfg[0]) );
    MUX2S_L muxa1(.o(da[1]),  .sel(f0), .i1(cfg[3]), .i0(cfg[2]) );
    MUX2S_L muxa2(.o(da[2]),  .sel(f0), .i1(cfg[5]), .i0(cfg[4]) );
    MUX2S_L muxa3(.o(da[3]),  .sel(f0), .i1(cfg[7]), .i0(cfg[6]) );
    MUX2S_L muxa4(.o(da[4]),  .sel(f0), .i1(cfg[9]), .i0(cfg[8]) );
    MUX2S_L muxa5(.o(da[5]),  .sel(f0), .i1(cfg[11]), .i0(cfg[10]) );
    MUX2S_L muxa6(.o(da[6]),  .sel(f0), .i1(cfg[13]), .i0(cfg[12]) );
    MUX2S_L muxa7(.o(da[7]),  .sel(f0), .i1(cfg[15]), .i0(cfg[14]) );
    MUX2S_L muxa8(.o(da[8]),  .sel(f0), .i1(cfg[17]), .i0(cfg[16]) );
    MUX2S_L muxa9(.o(da[9]),  .sel(f0), .i1(cfg[19]), .i0(cfg[18]) );
    MUX2S_L muxa10(.o(da[10]), .sel(f0), .i1(cfg[21]), .i0(cfg[20]) );
    MUX2S_L muxa11(.o(da[11]), .sel(f0), .i1(cfg[23]), .i0(cfg[22]) );
    MUX2S_L muxa12(.o(da[12]), .sel(f0), .i1(cfg[25]), .i0(cfg[24]) );
    MUX2S_L muxa13(.o(da[13]), .sel(f0), .i1(cfg[27]), .i0(cfg[26]) );
    MUX2S_L muxa14(.o(da[14]), .sel(f0), .i1(cfg[29]), .i0(cfg[28]) );
    MUX2S_L muxa15(.o(da[15]), .sel(f0), .i1(cfg[31]), .i0(cfg[30]) );

    MUX2S_L muxb0(.o(db[0]), .sel(f1), .i1(da[1]), .i0(da[0]) );
    MUX2S_L muxb1(.o(db[1]), .sel(f1), .i1(da[3]), .i0(da[2]) );
    MUX2S_L muxb2(.o(db[2]), .sel(f1), .i1(da[5]), .i0(da[4]) );
    MUX2S_L muxb3(.o(db[3]), .sel(f1), .i1(da[7]), .i0(da[6]) );
    MUX2S_L muxb4(.o(db[4]), .sel(f1), .i1(da[9]), .i0(da[8]) );
    MUX2S_L muxb5(.o(db[5]), .sel(f1), .i1(da[11]), .i0(da[10]) );
    MUX2S_L muxb6(.o(db[6]), .sel(f1), .i1(da[13]), .i0(da[12]) );
    MUX2S_L muxb7(.o(db[7]), .sel(f1), .i1(da[15]), .i0(da[14]) );

    MUX2S_L muxc0(.o(dc[0]), .sel(f2), .i1(db[1]), .i0(db[0]) );
    MUX2S_L muxc1(.o(dc[1]), .sel(f2), .i1(db[3]), .i0(db[2]) );
    MUX2S_L muxc2(.o(dc[2]), .sel(f2), .i1(db[5]), .i0(db[4]) );
    MUX2S_L muxc3(.o(dc[3]), .sel(f2), .i1(db[7]), .i0(db[6]) );

    MUX2S_L muxd0(.o(dd[0]), .sel(f3), .i1(dc[1]), .i0(dc[0]) );
    MUX2S_L muxd1(.o(dd[1]), .sel(f3), .i1(dc[3]), .i0(dc[2]) );

    MUX2S_L muxe0(.o(de), .sel(f4), .i1(dd[1]), .i0(dd[0]) );

    assign      dx = de;

	specify
       
	( f0 =>  dx    ) = (0,0);
	( f1 =>  dx    ) = (0,0);
	( f2 =>  dx    ) = (0,0);
	( f3 =>  dx    ) = (0,0);
	( f4 =>  dx    ) = (0,0);
	
     endspecify

`endif

endmodule

`endif
module MUX2S_L (
        o,
        sel,
        i0,
        i1
);

input        i0;
input        i1;
input        sel;

output        o;

`ifndef CS_SW_SKEL
	assign         o = (sel == 1'b0) ? i0 :
                    (sel == 1'b1) ? i1 :
                    (i0  == i1  ) ? i0 :1'bx;
    specify
        ( i0 =>  o ) = (0,0);
        ( i1 =>  o ) = (0,0);
        ( sel =>  o ) = (0,0);
    endspecify

`endif

endmodule
module OENC (
	f_oen,
	clk,
	gbl_clear_b,
	init_b,
	oen,
	rst,
	set_,
	CFG_OEN_INV,
	CFG_OEN_INV_,
	CFG_OEN_SEL
	);
output	f_oen;
input	clk,gbl_clear_b,init_b,oen,rst,set_;
input	CFG_OEN_INV;
input	CFG_OEN_INV_;
input	[3:0]	CFG_OEN_SEL;

wire	oen_inv;
assign oen_inv =({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b011) ? ~oen : 
				({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b101) ? oen :
				({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b000) ? 1'b0 :
				({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b001) ? 1'b0 : 1'bx;
reg		oen_psync;
reg		oen_nsync;

always @(posedge clk or posedge rst or negedge set_)
	if(~set_) oen_psync <= 1;
	else if(rst) oen_psync <= 0;
	else oen_psync <= oen_inv;
always @(negedge clk or posedge rst or negedge set_)
	if(~set_) oen_nsync <= 1;
	else if(rst) oen_nsync <= 0;
	else oen_nsync <= oen_inv;

wire	oen_sel;
assign oen_sel =({CFG_OEN_SEL,init_b} == 5'b00011) ? oen_nsync :
				({CFG_OEN_SEL,init_b} == 5'b00101) ? oen_psync :
				({CFG_OEN_SEL,init_b} == 5'b01001) ? oen_inv:
				({CFG_OEN_SEL,init_b} == 5'b10001) ? 1'b0:
				({CFG_OEN_SEL,init_b} == 5'b00000) ? 1'b1:
				({CFG_OEN_SEL,init_b} == 5'b00001) ? 1'b1 : 1'bx;
assign f_oen = !(gbl_clear_b & ~oen_sel);
endmodule


module co_lock_gate( TE, E, CP, Q);
input  TE;
input  E;
input  CP;
output Q;

wire en_t = E | TE;

reg en_latch;
always @(*) begin
    if (CP == 0)
        en_latch <= en_t;
end

assign Q = CP & en_latch;
endmodule

//Verilog HDL for "QC150_PLL_sim", "PLL_TOP" "functional"
`timescale 1ns/1ps

module PLL_TOP(
                 VDDIO        ,  //io power supply for regulator  
                 VSSIO        ,  //io ground for regulator
                 DVDD         ,  //digital power supply
                 DVSS         ,  //digital ground
                 AVSS_VCO     ,  //VCO ground
                 AVSS         ,  //analog ground
                 VREF         ,  //reference voltage for regulator
                 PDB          ,  //power-down mode control
                 RSTPLL       ,  //reset PLL control  
                 PLLCK0       ,  //PLL reference clock0
                 PLLCK1       ,  //PLL reference clock1
                 FBIN         ,  //feedback clock for deskew mode
                 CKSEL        ,  //PLL reference clk sel when ck_switch off
                 CK_SWITCH_EN ,  // Input clock automatic selection enable 0:manual select  (default) 1:automatic select
                 SEL_FBPATH   ,  //select the feedback signal to PFD  
                 DIVN         ,  //input divider control
                 DIVM         ,  //loop divider control
                 DIVFB        ,  //internal feedback clock of VCO control
                 LPF          ,  //loop filter resistance value adjustment
                 CPSEL_CR     ,  //select CP current,coarse tune
                 CPSEL_FN     ,  //select CP current,fine tune
                 CP_AUTO_ENB  ,  //cp current control sel
                 RST_REG_ENB  ,  //internal regulator por signal control
                 CALIB_EN     ,  // vco calibration enable 
                 CALIB_RSTN   ,  // vco calibration reset
                 CALIB_MANUAL ,  // vco calibration manual mode
                 CALIB_WIN    ,  // vco calibration vc monitor voltage window sel
                 CALIB_DIV    ,  // vco calibration manual mode
                 CALIB_16_32U ,  // vco calibration manual mode
                 BP_VDOUT     ,  //bypass dvdd(core) to vddd
                 LKD_MUX      ,  //lock detector ref clk sel 0: feedback clk 1:reference clk
                 FORCE_LOCK   ,  //force PLOCK signal to high
                 FLDD         ,  //lock detector range select
                 ATEST_EN     ,  //test control enable for analog test 
                 DTEST_EN     ,  //test control enable for digital test 
                 ATEST_SEL    ,  //analog test select
                 DTEST_SEL    ,  //digital test select
                 VCO_INI_SEL  ,  //vco initial phase align control
                 LKD_TOL      ,  //Lock Detector tolerance (TBD)
                 LKD_HOLD     ,  // Lock Detector hold number (TBD) 
                 VRSEL        ,  //select the reference voltage for regulator
                 BK           ,  //Back up register 
                 SSEN         ,  //Spread spectrum function enable 0:don't use SSCG function  (default) 1:enable
                 SSDIVH       ,  //Spread frequency-divider 1 control, range within[1,16] divider value NH=SSDIVH<3:0>+1
                 SSDIVL       ,  //Spread frequency-divider 2 control, range within[1,256] divider value NH=SSDIVL<7:0>+1
                 SSRG         ,  //Spread ratio select (TBD)
                 PSEN         ,  // dynamic phase shift enable
                 PSCK         ,  // dynamic phase shift clock
                 PSDIR        ,  // dynamic phase shift direction
                 PSSEL        ,  // dynamic phase shift channel sel                 
                 MKEN0        ,  //output enable for channel 0
                 MKEN1        ,  //output enable for channel 1
                 MKEN2        ,  //output enable for channel 2
                 MKEN3        ,  //output enable for channel 3
                 MKEN4        ,  //output enable for channel 4
                 MKEN5        ,  //output enable for channel 5
                 BPS0         ,  //bypass output of channel 0
                 BPS1         ,  //bypass output of channel 1
                 BPS2         ,  //bypass output of channel 2
                 BPS3         ,  //bypass output of channel 3
                 BPS4         ,  //bypass output of channel 4
                 BPS5         ,  //bypass output of channel 5
                 FRAC         ,  //Frac-divider setting
                 DIVC0        ,  //output divider control for channel 0
                 DIVC1        ,  //output divider control for channel 1
                 DIVC2        ,  //output divider control for channel 2
                 DIVC3        ,  //output divider control for channel 3
                 DIVC4        ,  //output divider control for channel 4
                 DIVC5        ,  //output divider control for channel 5
                 CO0DLY       ,  //channel 0 coarse delay control
                 CO1DLY       ,  //channel 1 coarse delay control
                 CO2DLY       ,  //channel 2 coarse delay control
                 CO3DLY       ,  //channel 3 coarse delay control
                 CO4DLY       ,  //channel 4 coarse delay control
                 CO5DLY       ,  //channel 5 coarse delay control
                 P0SEL        ,  //select phase for channel 0
                 P1SEL        ,  //select phase for channel 1
                 P2SEL        ,  //select phase for channel 2
                 P3SEL        ,  //select phase for channel 3
                 P4SEL        ,  //select phase for channel 4
                 P5SEL        ,  //select phase for channel 5
                 PFBSEL       ,  //select phase for CKFB
                 CO0          ,  //PLL output clock channel 0
                 CO1          ,  //PLL output clock channel 1
                 CO2          ,  //PLL output clock channel 2
                 CO3          ,  //PLL output clock channel 3
                 CO4          ,  //PLL output clock channel 4
                 CO5          ,  //PLL output clock channel 5
                 FBOUT        ,  //PLL feedback clock
                 ACTIVECK     ,  //Indicated that which clock is selected now
                 CKBAD0       ,  //Indicated PLLCK0 clock is bad
                 CKBAD1       ,  //Indicated PLLCK1 clock is bad
                 PSDONE       ,  // dynamic phase shift status flag
                 PLOCK        ,  //PLL lock status output
                 ATEST_PLL    ,  //analog signal test output
                 DTEST_PLL       //digital signal test output                           
             );

//port definition

input         VDDIO        ;  //io power supply for regulator  
input         VSSIO        ;  //io ground for regulator
input         DVDD         ;  //digital power supply
input         DVSS         ;  //digital ground
input         AVSS_VCO     ;  //VCO ground
input         AVSS         ;  //analog ground
input         PLLCK0       ;  //PLL reference clock0
input         PLLCK1       ;  //PLL reference clock1
input         FBIN         ;  //feedback clock for deskew mode
input         VREF         ;  //reference voltage for regulator
input         CKSEL        ;  //PLL reference clk sel when ck_switch off
input         CK_SWITCH_EN ;  // Input clock automatic selection enable 0:manual select  (default) 1:automatic select
input         PDB          ;  //power-down mode control
input         RSTPLL       ;  //reset PLL control
input         SEL_FBPATH   ;  //select the feedback signal to PFD

input  [7:0]  DIVN         ;  //input divider control
input  [7:0]  DIVM         ;  //loop divider control
input         DIVFB        ;  //internal feedback clock of VCO control 1:bypass. 0:divide by 2

input  [2:0]  LPF          ;  //loop filter resistance value adjustment
input  [2:0]  CPSEL_CR     ;  //select CP current,coarse tune
input  [6:0]  CPSEL_FN     ;  //select CP current,fine tune
input         CP_AUTO_ENB  ;  //cp current control sel
input         RST_REG_ENB  ;  //internal regulator por signal control
input         CALIB_EN     ;  // vco calibration enable 
input         CALIB_RSTN   ;  // vco calibration reset
input  [3:0]  CALIB_MANUAL ;  // vco calibration manual mode
input  [1:0]  CALIB_WIN    ;  // vco calibration vc monitor voltage window sel
input  [7:0]  CALIB_DIV    ;  // vco calibration clock divider setting
input         CALIB_16_32U ;  // vco calibration time sel
input         BP_VDOUT     ;  //bypass dvdd(core) to vddd
input         LKD_MUX      ;  //lock detector ref clk sel 0: feedback clk 1:reference clk
input         FORCE_LOCK   ;  //force PLOCK signal to high
input  [1:0]  FLDD         ;  //lock detector range select
input         ATEST_EN     ;  //test control enable for analog test 
input         DTEST_EN     ;  //test control enable for digital test 
input         ATEST_SEL    ;  //analog test select
input         DTEST_SEL    ;  //digital test select
input         VCO_INI_SEL  ;  //vco initial phase align control
input         LKD_TOL      ;  //Lock Detector tolerance (TBD)
input         LKD_HOLD     ;  // Lock Detector hold number (TBD) 
input  [1:0]  VRSEL        ;  //select the reference voltage for regulator
input  [3:0]  BK           ;  //Back up register 

input         SSEN         ;  //Spread spectrum function enable 0:don't use SSCG function  (default) 1:enable
input  [1:0]  SSDIVH       ;  //Spread frequency-divider 1 control, range within[1,16] divider value NH=SSDIVH<3:0>+1
input  [7:0]  SSDIVL       ;  //Spread frequency-divider 2 control, range within[1,256] divider value NH=SSDIVL<7:0>+1
input  [1:0]  SSRG         ;  //Spread ratio select (TBD)
input         PSEN         ;  // dynamic phase shift enable
input         PSCK         ;  // dynamic phase shift clock
input         PSDIR        ;  // dynamic phase shift direction
input  [5:0]  PSSEL        ;  // dynamic phase shift channel sel

input         MKEN0        ;  //output enable for channel 0
input         MKEN1        ;  //output enable for channel 1
input         MKEN2        ;  //output enable for channel 2
input         MKEN3        ;  //output enable for channel 3
input         MKEN4        ;  //output enable for channel 4
input         MKEN5        ;  //output enable for channel 5
input         BPS0         ;  //bypass output of channel 0
input         BPS1         ;  //bypass output of channel 1
input         BPS2         ;  //bypass output of channel 2
input         BPS3         ;  //bypass output of channel 3
input         BPS4         ;  //bypass output of channel 4
input         BPS5         ;  //bypass output of channel 5
input  [2:0]  FRAC         ;  //Frac-divider setting
input  [7:0]  DIVC0        ;  //output divider control for channel 0
input  [7:0]  DIVC1        ;  //output divider control for channel 1
input  [7:0]  DIVC2        ;  //output divider control for channel 2
input  [7:0]  DIVC3        ;  //output divider control for channel 3
input  [7:0]  DIVC4        ;  //output divider control for channel 4
input  [7:0]  DIVC5        ;  //output divider control for channel 5
input  [7:0]  CO0DLY       ;  //channel 0 coarse delay control
input  [7:0]  CO1DLY       ;  //channel 1 coarse delay control
input  [7:0]  CO2DLY       ;  //channel 2 coarse delay control
input  [7:0]  CO3DLY       ;  //channel 3 coarse delay control
input  [7:0]  CO4DLY       ;  //channel 4 coarse delay control
input  [7:0]  CO5DLY       ;  //channel 5 coarse delay control
input  [2:0]  P0SEL        ;  //select phase for channel 0
input  [2:0]  P1SEL        ;  //select phase for channel 1
input  [2:0]  P2SEL        ;  //select phase for channel 2
input  [2:0]  P3SEL        ;  //select phase for channel 3
input  [2:0]  P4SEL        ;  //select phase for channel 4
input  [2:0]  P5SEL        ;  //select phase for channel 5
input  [2:0]  PFBSEL       ;  //select phase for feedback clock

output        CO0          ;  //PLL output clock channel 0
output        CO1          ;  //PLL output clock channel 1
output        CO2          ;  //PLL output clock channel 2
output        CO3          ;  //PLL output clock channel 3
output        CO4          ;  //PLL output clock channel 4
output        CO5          ;  //PLL output clock channel 5
output        FBOUT        ;  //PLL feedback clock output
output        ACTIVECK     ;  //Indicated that which clock is selected now
output        CKBAD0       ;  //Indicated PLLCK0 clock is bad
output        CKBAD1       ;  //Indicated PLLCK1 clock is bad
output        PSDONE       ;  // dynamic phase shift status flag
output        PLOCK        ;  //PLL lock status output
output        ATEST_PLL    ;  //analog signal test output
output        DTEST_PLL    ;  //digital signal test output


//parameters definition

parameter MAX_INPUT_PERIOD   = 100;    // input freq       : 10MHZ--700MHz
parameter MIN_INPUT_PERIOD   = 1.428;         //
parameter MAX_PFD_PERIOD     = 100;        // PFD input freq   : 10MHZ--450MHz
parameter MIN_PFD_PERIOD     = 2.222;          //
parameter MAX_VCO_PERIOD     = 1.667;        // VCO operate freq : 600MHZ--1400MHz
parameter MIN_VCO_PERIOD     = 0.714;          //
parameter MAX_OUTPUT_PERIOD  = 854.7;        // output freq      : 1.17MHZ--700MHz
parameter MIN_OUTPUT_PERIOD  = 1.428;          //
parameter LOCK_TIME          = 10;       //lock time range is several us. Now we set the default value 10ps.

//internal signal definition
wire  ck_bps;
wire  refck;
wire  ckin;
wire  fs_input_range;
wire  fs_pfd_range;
wire  fs_vco_range;
wire  dsk_input_range;
wire  dsk_pfd_range;
wire  dsk_vco_range;
wire  lock_pd;
wire  lock_fl;
wire  lock_fs;
wire  lock_dsk;
wire  lock_val_loop;
wire  lock_val;
wire  [5:0]  lock_th;
reg   [5:0]  lock_cnt;
reg   lock_tmp;
reg   PLOCK;
reg   plock_en;
wire  [8:0]  divn_num;
wire  [8:0]  divm_num;
wire  [1:0]  divfb_num;
wire  [2:0]  frac_num;
wire  [8:0]  divc0_num;
wire  [8:0]  divc1_num;
wire  [8:0]  divc2_num;
wire  [8:0]  divc3_num;
wire  [8:0]  divc4_num;
wire  [8:0]  divc5_num;
wire  [8:0]  divcfb_num;
reg   vco_mp_tmp;
reg   [7:0]  vco_mp_p;
wire  vco_mp_loop;

wire  C0_sel;
wire  C0_rb_en;
wire  C0_rb;
reg   C0_clk_tmp;
reg   C0_rb_tmp;
reg   [7:0]  C0_dlycnt;
wire  C0_divcnt_en;
reg   C0_phase_align;
wire  C0_out_tmp;

wire  C1_sel;
wire  C1_rb_en;
wire  C1_rb;
reg   C1_clk_tmp;
reg   C1_rb_tmp;
reg   [7:0]  C1_dlycnt;
wire  C1_divcnt_en;
reg   C1_phase_align;
wire  C1_out_tmp;

wire  C2_sel;
wire  C2_rb_en;
wire  C2_rb;
reg   C2_clk_tmp;
reg   C2_rb_tmp;
reg   [7:0]  C2_dlycnt;
wire  C2_divcnt_en;
reg   C2_phase_align;
wire  C2_out_tmp;

wire  C3_sel;
wire  C3_rb_en;
wire  C3_rb;
reg   C3_clk_tmp;
reg   C3_rb_tmp;
reg   [7:0]  C3_dlycnt;
wire  C3_divcnt_en;
reg   C3_phase_align;
wire  C3_out_tmp;

wire  C4_sel;
wire  C4_rb_en;
wire  C4_rb;
reg   C4_clk_tmp;
reg   C4_rb_tmp;
reg   [7:0]  C4_dlycnt;
wire  C4_divcnt_en;
reg   C4_phase_align;
wire  C4_out_tmp;

wire  C5_sel;
wire  C5_rb_en;
wire  C5_rb;
reg   C5_clk_tmp;
reg   C5_rb_tmp;
reg   [7:0]  C5_dlycnt;
wire  C5_divcnt_en;
reg   C5_phase_align;
wire  C5_out_tmp;

wire  CFB_sel;
wire  CFB_rb_en;
wire  CFB_rb;
reg   CFB_clk_tmp;
reg   CFB_rb_tmp;
reg   [7:0]  CFB_dlycnt;
wire  CFB_divcnt_en;
reg   CFB_phase_align;
wire  CFB_out_tmp;


realtime t1;
realtime t2;
real  period_in; //integer period_in;
real  period_mp; //integer period_mp;
real  divc0_frac;
real  period_c0;
real  period_c1;
real  period_c2;
real  period_c3;
real  period_c4;
real  period_c5;
real  period_cFB;

//initial the state

  initial begin
        period_in  = 50.000;
        period_mp  = 50.000;
        t1         = 50;
        t2         = 0;

  end

  assign lock_th = 6'b111111;
  assign divn_num = DIVN + 9'd1;
  assign divm_num = DIVM + 9'd1;
  assign divfb_num = DIVFB + 1'b1;
  
  assign divc0_num = DIVC0 + 9'd1;
  assign frac_num  = FRAC;  
  assign divc1_num = DIVC1 + 9'd1;
  assign divc2_num = DIVC2 + 9'd1;
  assign divc3_num = DIVC3 + 9'd1;
  assign divc4_num = DIVC4 + 9'd1;
  assign divc5_num = DIVC5 + 9'd1;
  
//detect the input clock period


 assign refck = (CKSEL == 0 ) ? PLLCK0 : PLLCK1;

 assign ckin = (PDB==1'b0 || refck == 1'bz || refck == 1'bx) ? 1'b0 : refck;
                                                               
 assign ck_bps = (refck == 1'bz || refck == 1'bx) ? 1'b0 : refck;

 always @(posedge ckin) begin
        
        t2  = t2- t1 > 1000 
            ? $realtime - 50
            : t1 - t2 > 1000
              ? $realtime - 50
              : t1;
        t1=$realtime;


        if(t2 == 50) 
          period_in = 50;
        else if (t1-t2 > 210 || t2-t1 > 210 || period_in > 210)
          period_in = 210;
        else if (period_in < 5)
          period_in = 5;
        else
          period_in = t1 -t2;
 end

//lock judgement

  assign fs_input_range = ((period_in <= MAX_INPUT_PERIOD) && (period_in >= MIN_INPUT_PERIOD)) ? 1'b1 : 1'b0;
  assign fs_pfd_range = ((period_in*divn_num <= MAX_PFD_PERIOD) && (period_in*divn_num >= MIN_PFD_PERIOD)) ? 1'b1 : 1'b0;
  assign fs_vco_range = ((period_in*divn_num/(divm_num*divfb_num) <= MAX_VCO_PERIOD) && (period_in*divn_num/(divm_num*divfb_num) >= MIN_VCO_PERIOD)) ? 1'b1 : 1'b0;
  assign dsk_input_range = ((period_in <= MAX_INPUT_PERIOD) && (period_in >= MIN_INPUT_PERIOD)) ? 1'b1 : 1'b0;
  assign dsk_pfd_range = ((period_in*divn_num <= MAX_PFD_PERIOD) && (period_in*divn_num >= MIN_PFD_PERIOD)) ? 1'b1 : 1'b0;
  assign dsk_vco_range = ((period_in*divn_num/(divm_num*divfb_num) <= MAX_VCO_PERIOD) && (period_in*divn_num/(divm_num*divfb_num) >= MIN_VCO_PERIOD)) ? 1'b1 : 1'b0;
  assign lock_pd = 1'b0;
  assign lock_fl = 1'b1;
  assign lock_fs = (fs_input_range && fs_pfd_range && fs_vco_range) ? 1'b1 : 1'b0;
  assign lock_dsk = (dsk_input_range && dsk_pfd_range && dsk_vco_range) ? 1'b1 : 1'b0;
  assign lock_val_loop = (RSTPLL || !PDB) ? lock_pd :
        (!SEL_FBPATH) ? lock_fs : lock_dsk ;
  assign lock_val = (RSTPLL || !PDB) ? lock_pd :
                    FORCE_LOCK ? lock_fl : lock_val_loop;
  initial begin
  lock_cnt = 6'b000000;
  lock_tmp = 1'b0;
  PLOCK = 1'b0;
  end 
  always @(posedge ckin) begin
  if (lock_val == 1'b0) begin
        lock_tmp <= 1'b0;
        lock_cnt <= 6'b000000;
            end
  else if (lock_cnt[5:0] == lock_th[5:0]) begin
         lock_tmp <= 1'b1;
         lock_cnt <= lock_th[5:0];
                end
  else lock_cnt <= lock_cnt + 7'd1;
  end

  always @(posedge lock_tmp) PLOCK <= #LOCK_TIME lock_tmp;
  always @(negedge lock_tmp) PLOCK <= lock_tmp;

//PLL loop model

  initial begin
  vco_mp_tmp = 1'b0;
  vco_mp_p = 8'b00000000;
  end

  always @(SEL_FBPATH  or period_in or divn_num or divm_num or divfb_num) begin
  if (!SEL_FBPATH) period_mp = period_in*divn_num/(divm_num*divfb_num*1.000);
  else             period_mp = period_in*divn_num/(divm_num*divfb_num*1.000);
  end

 
  initial begin
    wait (VDDIO);
    #300;
    forever vco_mp_tmp = #(period_mp/2.000) !vco_mp_tmp;
    
  end

  assign vco_mp_loop = (!PDB || RSTPLL) ? 1'b0 :
      (lock_val_loop) ? vco_mp_tmp : 1'b0;
  always @(negedge vco_mp_loop or negedge PDB or posedge RSTPLL) 
  if (!PDB || RSTPLL) plock_en <= 1'b0;
  else        plock_en <= PLOCK;
  
 always @(plock_en or vco_mp_loop or period_mp) begin
  if (!plock_en) vco_mp_p = 8'b00000000;
  else begin  vco_mp_p[0] <= vco_mp_loop;
      vco_mp_p[1] <= #(1*period_mp/8.000) vco_mp_loop;  
      vco_mp_p[2] <= #(2*period_mp/8.000) vco_mp_loop;  
      vco_mp_p[3] <= #(3*period_mp/8.000) vco_mp_loop;  
      vco_mp_p[4] <= #(4*period_mp/8.000) vco_mp_loop;  
      vco_mp_p[5] <= #(5*period_mp/8.000) vco_mp_loop;  
      vco_mp_p[6] <= #(6*period_mp/8.000) vco_mp_loop;  
      vco_mp_p[7] <= #(7*period_mp/8.000) vco_mp_loop;
       end  
  end

//output C0 assignment

  assign C0_sel = (P0SEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (P0SEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (P0SEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (P0SEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (P0SEL[2:0] == 3'b100) ? vco_mp_p[4] :
      (P0SEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (P0SEL[2:0] == 3'b110) ? vco_mp_p[6] :
                               vco_mp_p[7] ;

  always @(frac_num or divc0_frac or divc0_num) begin
        
   divc0_frac = frac_num*0.125 + divc0_num;
        
  end

  assign C0_rb_en = (PDB && !RSTPLL && MKEN0) ? 1'b1 : 1'b0;
  assign C0_rb = (PLOCK && C0_rb_en) ? 1'b1 : 1'b0;
  always @(negedge C0_sel or negedge C0_rb) begin
  if (!C0_rb)  C0_rb_tmp <= 1'b0;
  else    C0_rb_tmp <= 1'b1;
  end
  always @(posedge C0_sel or negedge C0_rb_tmp) begin
  if (!C0_rb_tmp)        C0_dlycnt <= 8'd0;
  else if (C0_dlycnt[7:0] == CO0DLY[7:0] + 8'd1)  C0_dlycnt <= CO0DLY[7:0] + 8'd1;
  else          C0_dlycnt <= C0_dlycnt + 8'd1;
  end

  assign C0_divcnt_en = (C0_dlycnt[7:0] == CO0DLY[7:0]  + 8'd1); 
  
  always @(period_mp or divc0_frac) begin

     period_c0 = period_mp*divc0_frac;

  end

  initial begin
  C0_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    C0_phase_align  <= 1'b0;
    C0_clk_tmp      <= 1'b0;
    wait (C0_phase_align);
    forever   C0_clk_tmp = #(period_c0/2.000) !C0_clk_tmp;
   
  end
  

  always @(posedge C0_sel) begin

    if (C0_divcnt_en && C0_rb_tmp)  C0_phase_align  <= 1'b1;
  
  end

   
  assign C0_out_tmp = C0_clk_tmp;


  assign CO0 = (BPS0) ? ck_bps : C0_out_tmp ;

//output C1 assignment

assign C1_sel = (P1SEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (P1SEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (P1SEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (P1SEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (P1SEL[2:0] == 3'b100) ? vco_mp_p[4] :
      (P1SEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (P1SEL[2:0] == 3'b110) ? vco_mp_p[6] :
                     vco_mp_p[7] ;
  assign C1_rb_en = (PDB && !RSTPLL && MKEN1) ? 1'b1 : 1'b0;
  assign C1_rb = (PLOCK && C1_rb_en) ? 1'b1 : 1'b0;
  always @(negedge C1_sel or negedge C1_rb) begin
  if (!C1_rb)  C1_rb_tmp <= 1'b0;
  else    C1_rb_tmp <= 1'b1;
  end
  always @(posedge C1_sel or negedge C1_rb_tmp) begin
  if (!C1_rb_tmp)        C1_dlycnt <= 8'd0;
  else if (C1_dlycnt[7:0] == CO1DLY[7:0] + 8'd1 )  C1_dlycnt <= CO1DLY[7:0] + 8'd1 ;
  else          C1_dlycnt <= C1_dlycnt + 8'd1;
  end

  assign C1_divcnt_en = (C1_dlycnt[7:0] == CO1DLY[7:0] + 8'd1) ;
  
  always @(period_mp or divc1_num) begin

     period_c1 = period_mp*divc1_num;

  end

  initial begin
  C1_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    C1_phase_align  <= 1'b0;
    C1_clk_tmp      <= 1'b0;
    wait (C1_phase_align);
    forever   C1_clk_tmp = #(period_c1/2.000) !C1_clk_tmp;
   
  end
  

  always @(posedge C1_sel) begin

    if (C1_divcnt_en && C1_rb_tmp)  C1_phase_align  <= 1'b1;
  
  end

   
  assign C1_out_tmp = C1_clk_tmp;

   
  assign CO1 = (BPS1) ? ck_bps : C1_out_tmp ;
 
//output C2 assignment

assign C2_sel = (P2SEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (P2SEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (P2SEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (P2SEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (P2SEL[2:0] == 3'b100) ? vco_mp_p[4] :
      (P2SEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (P2SEL[2:0] == 3'b110) ? vco_mp_p[6] :
                     vco_mp_p[7] ;
  assign C2_rb_en = (PDB && !RSTPLL && MKEN2) ? 1'b1 : 1'b0;
  assign C2_rb = (PLOCK && C2_rb_en) ? 1'b1 : 1'b0;
  always @(negedge C2_sel or negedge C2_rb) begin
  if (!C2_rb)  C2_rb_tmp <= 1'b0;
  else    C2_rb_tmp <= 1'b1;
  end
  always @(posedge C2_sel or negedge C2_rb_tmp) begin
  if (!C2_rb_tmp)        C2_dlycnt <= 8'd0;
  else if (C2_dlycnt[7:0] == CO2DLY[7:0] + 8'd1 )  C2_dlycnt <= CO2DLY[7:0] + 8'd1 ;
  else          C2_dlycnt <= C2_dlycnt + 8'd1;
  end

  assign C2_divcnt_en = (C2_dlycnt[7:0] == CO2DLY[7:0] + 8'd1) ;
  
  always @(period_mp or divc2_num) begin

     period_c2 = period_mp*divc2_num;

  end

  initial begin
  C2_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    C2_phase_align  <= 1'b0;
    C2_clk_tmp      <= 1'b0;
    wait (C2_phase_align);
    forever   C2_clk_tmp = #(period_c2/2.000) !C2_clk_tmp;
   
  end
  

  always @(posedge C2_sel) begin

    if (C2_divcnt_en && C2_rb_tmp)  C2_phase_align  <= 1'b1;
  
  end

   
  assign C2_out_tmp = C2_clk_tmp;

   
  assign CO2 = (BPS2) ? ck_bps : C2_out_tmp ;
 
//output C3 assignment

assign C3_sel = (P3SEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (P3SEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (P3SEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (P3SEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (P3SEL[2:0] == 3'b100) ? vco_mp_p[4] :
      (P3SEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (P3SEL[2:0] == 3'b110) ? vco_mp_p[6] :
                     vco_mp_p[7] ;
  assign C3_rb_en = (PDB && !RSTPLL && MKEN3) ? 1'b1 : 1'b0;
  assign C3_rb = (PLOCK && C3_rb_en) ? 1'b1 : 1'b0;
  always @(negedge C3_sel or negedge C3_rb) begin
  if (!C3_rb)  C3_rb_tmp <= 1'b0;
  else    C3_rb_tmp <= 1'b1;
  end
  always @(posedge C3_sel or negedge C3_rb_tmp) begin
  if (!C3_rb_tmp)        C3_dlycnt <= 8'd0;
  else if (C3_dlycnt[7:0] == CO3DLY[7:0] + 8'd1 )  C3_dlycnt <= CO3DLY[7:0] + 8'd1 ;
  else          C3_dlycnt <= C3_dlycnt + 8'd1;
  end

  assign C3_divcnt_en = (C3_dlycnt[7:0] == CO3DLY[7:0] + 8'd1) ;
  
  always @(period_mp or divc3_num) begin

     period_c3 = period_mp*divc3_num;

  end

  initial begin
  C3_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    C3_phase_align  <= 1'b0;
    C3_clk_tmp      <= 1'b0;
    wait (C3_phase_align);
    forever   C3_clk_tmp = #(period_c3/2.000) !C3_clk_tmp;
   
  end
  

  always @(posedge C3_sel) begin

    if (C3_divcnt_en && C3_rb_tmp)  C3_phase_align  <= 1'b1;
  
  end

   
  assign C3_out_tmp = C3_clk_tmp;

   
  assign CO3 = (BPS3) ? ck_bps : C3_out_tmp ;

//output C4 assignment

assign C4_sel = (P4SEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (P4SEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (P4SEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (P4SEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (P4SEL[2:0] == 3'b100) ? vco_mp_p[4] :
      (P4SEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (P4SEL[2:0] == 3'b110) ? vco_mp_p[6] :
                     vco_mp_p[7] ;
  assign C4_rb_en = (PDB && !RSTPLL && MKEN4) ? 1'b1 : 1'b0;
  assign C4_rb = (PLOCK && C4_rb_en) ? 1'b1 : 1'b0;
  always @(negedge C4_sel or negedge C4_rb) begin
  if (!C4_rb)  C4_rb_tmp <= 1'b0;
  else    C4_rb_tmp <= 1'b1;
  end
  always @(posedge C4_sel or negedge C4_rb_tmp) begin
  if (!C4_rb_tmp)        C4_dlycnt <= 8'd0;
  else if (C4_dlycnt[7:0] == CO4DLY[7:0] + 8'd1 )  C4_dlycnt <= CO4DLY[7:0] + 8'd1 ;
  else          C4_dlycnt <= C4_dlycnt + 8'd1;
  end

  assign C4_divcnt_en = (C4_dlycnt[7:0] == CO4DLY[7:0] + 8'd1) ;
  
  always @(period_mp or divc4_num) begin

     period_c4 = period_mp*divc4_num;

  end

  initial begin
  C4_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    C4_phase_align  <= 1'b0;
    C4_clk_tmp      <= 1'b0;
    wait (C4_phase_align);
    forever   C4_clk_tmp = #(period_c4/2.000) !C4_clk_tmp;
   
  end
  

  always @(posedge C4_sel) begin

    if (C4_divcnt_en && C4_rb_tmp)  C4_phase_align  <= 1'b1;
  
  end

   
  assign C4_out_tmp = C4_clk_tmp;

   
  assign CO4 = (BPS4) ? ck_bps : C4_out_tmp ;

//output C5 assignment

assign C5_sel = (P5SEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (P5SEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (P5SEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (P5SEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (P5SEL[2:0] == 3'b100) ? vco_mp_p[5] :
      (P5SEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (P5SEL[2:0] == 3'b110) ? vco_mp_p[6] :
                     vco_mp_p[7] ;
  assign C5_rb_en = (PDB && !RSTPLL && MKEN5) ? 1'b1 : 1'b0;
  assign C5_rb = (PLOCK && C5_rb_en) ? 1'b1 : 1'b0;
  always @(negedge C5_sel or negedge C5_rb) begin
  if (!C5_rb)  C5_rb_tmp <= 1'b0;
  else    C5_rb_tmp <= 1'b1;
  end
  always @(posedge C5_sel or negedge C5_rb_tmp) begin
  if (!C5_rb_tmp)        C5_dlycnt <= 8'd0;
  else if (C5_dlycnt[7:0] == CO5DLY[7:0] + 8'd1 )  C5_dlycnt <= CO5DLY[7:0] + 8'd1 ;
  else          C5_dlycnt <= C5_dlycnt + 8'd1;
  end

  assign C5_divcnt_en = (C5_dlycnt[7:0] == CO5DLY[7:0] + 8'd1) ;
  
  always @(period_mp or divc5_num) begin

     period_c5 = period_mp*divc5_num;

  end

  initial begin
  C5_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    C5_phase_align  <= 1'b0;
    C5_clk_tmp      <= 1'b0;
    wait (C5_phase_align);
    forever   C5_clk_tmp = #(period_c5/2.000) !C5_clk_tmp;
   
  end
  

  always @(posedge C5_sel) begin

    if (C5_divcnt_en && C5_rb_tmp)  C5_phase_align  <= 1'b1;
  
  end

   
  assign C5_out_tmp = C5_clk_tmp;

   
  assign CO5 = (BPS5) ? ck_bps : C5_out_tmp ;

//output CFB assignment

assign CFB_sel = (PFBSEL[2:0] == 3'b000) ? vco_mp_p[0] :
      (PFBSEL[2:0] == 3'b001) ? vco_mp_p[1] :
      (PFBSEL[2:0] == 3'b010) ? vco_mp_p[2] :
      (PFBSEL[2:0] == 3'b011) ? vco_mp_p[3] :
      (PFBSEL[2:0] == 3'b100) ? vco_mp_p[4] :
      (PFBSEL[2:0] == 3'b101) ? vco_mp_p[5] :
      (PFBSEL[2:0] == 3'b110) ? vco_mp_p[6] :
                     vco_mp_p[7] ;
  assign CFB_rb_en = (PDB && !RSTPLL) ? 1'b1 : 1'b0;
  assign CFB_rb = ( CFB_rb_en) ? 1'b1 : 1'b0;
  always @(negedge CFB_sel or negedge CFB_rb) begin
  if (!CFB_rb)  CFB_rb_tmp <= 1'b0;
  else    CFB_rb_tmp <= 1'b1;
  end
  always @(posedge CFB_sel or negedge CFB_rb_tmp) begin
  if (!CFB_rb_tmp)        CFB_dlycnt <= 8'd0;
  else if (CFB_dlycnt[7:0] ==  8'd1 )  CFB_dlycnt <=  8'd1 ;
  else          CFB_dlycnt <= CFB_dlycnt + 8'd1;
  end

  assign CFB_divcnt_en = (CFB_dlycnt[7:0] ==  8'd1) ;
  
  always @(period_mp or divm_num) begin

     period_cFB = period_mp*divm_num;

  end

  initial begin
  CFB_clk_tmp = 1'b0;
  end
 
  initial begin
    wait (VDDIO);
    #300;
    CFB_phase_align  <= 1'b0;
    CFB_clk_tmp      <= 1'b0;
    wait (CFB_phase_align);
    forever   CFB_clk_tmp = #(period_cFB/2.000) !CFB_clk_tmp;
   
  end
  

  always @(posedge CFB_sel) begin

    if (CFB_divcnt_en && CFB_rb_tmp)  CFB_phase_align  <= 1'b1;
  
  end

   
  assign CFB_out_tmp = CFB_clk_tmp;

   
  assign FBOUT = CFB_out_tmp ;
 
endmodule



module CSGPIO (
     TXD
    ,TED
    ,RXD
    ,PAD
    ,NS_LV
    ,PDR
    ,NDR
    ,KEEP
    ,RX_DIG_EN
    ,VPCI_EN
);

input TXD;                    // data output to PDA
input TED;                    // data output enable
output RXD;                   // data input from PAD 
inout PAD;                    // PAD

// ------------- total 106 config bits
input [1:0] NS_LV;         // slew rate control
input [3:0] PDR;           // driving strength, P
input [3:0] NDR;           // driving strength, N
input [1:0] KEEP;          // pullup,pulldown,bus-keeper

input RX_DIG_EN;           // LVCMOS RX enable

input VPCI_EN;             // PCI diode enable
//--------------
 
supply1 VDDIO, VDDCORE;
supply0 VSSIO, VSSCORE;

    /* rx */

    wire rxe;
    
    assign rxe=~(RX_DIG_EN);
    bufif1 rx00 (RXD,PAD,RX_DIG_EN);
    nmos  NMOSrx0 (RXD, VSSIO, rxe);


    //------- driver 
//------LVCMOS  
    wire pdr0a,ndr0a,pdr0b,ndr0b,pdr0c,ndr0c,pdr1a,ndr1a,pdr1b,ndr1b,pdr1c,ndr1c;
      
    assign pdr0a=PDR[0]|PDR[1]|PDR[2]|PDR[3];
    assign ndr0a=NDR[0]|NDR[1]|NDR[2]|NDR[3];
    assign pdr0b=pdr0a&(NS_LV[0]|NS_LV[1])&(!TED);
    assign ndr0b=ndr0a&(NS_LV[0]|NS_LV[1])&(!TED);
    assign pdr0c=~( pdr0b & TXD );
    assign ndr0c=~(!ndr0b | TXD );
    
    pmos  pdriver00 (PAD, VDDIO, pdr0c);
    nmos  ndriver00 (PAD, VSSIO, ndr0c);


    
    //--------- Pullup 
    wire pullup0,pullup1,pulldn0,pulldn1;
    
    assign pullup0=~(KEEP[1]&((!KEEP[0])|(KEEP[0]&!RXD)));
    
    rpmos    PMOS0A    (PAD,        PAD0PA_out, pullup0);
    rpmos    PMOS0B    (PAD0PA_out, PAD0PB_out, pullup0);
    rpmos    PMOS0C    (PAD0PB_out, VDDIO,      pullup0);    


    //---------- Pulldown (Strength to Weak)
    assign pulldn0=(KEEP[0]&((!KEEP[1])|(KEEP[1]&RXD)));
    
    rnmos    NMOS0A    (PAD,        PAD0NA_out, pulldn0);
    rnmos    NMOS0B    (PAD0NA_out, PAD0NB_out, pulldn0);
    rnmos    NMOS0C    (PAD0NB_out, VSSIO,      pulldn0);

    
    //-------- keeper 

endmodule

module io_data(
     f_oen
    ,f_od
    ,id
    ,ted
    ,txd
    ,rxd
    ,CFG_OEN_SEL
    ,CFG_OUT_SEL
);

input          f_oen;
input          f_od;
output         id;
output         ted;
output         txd;
input          rxd;
input  [1:0]   CFG_OEN_SEL;
input  [1:0]   CFG_OUT_SEL;

assign ted = CFG_OEN_SEL == 2'b00 ?  1'b1  :
             CFG_OEN_SEL == 2'b01 ?  1'b0  :
             CFG_OEN_SEL == 2'b10 ?  f_oen :
             CFG_OEN_SEL == 2'b11 ? ~f_oen :
                                     1'bx  ;

assign txd = CFG_OUT_SEL == 2'b00 ?  1'b1  :
             CFG_OUT_SEL == 2'b01 ?  1'b0  :
             CFG_OUT_SEL == 2'b10 ?  f_od  :
             CFG_OUT_SEL == 2'b11 ? ~f_od  :
                                     1'bx  ;
assign id = rxd;

endmodule

//MUX2S1 & iob_dff used in UPDATE module
module IO_MUX2S1(
	o,
	in0,
	in1,
	SEL
	);
output	o;
input	in0;
input	in1;
input	SEL;

assign o = SEL ? in1 : in0;
endmodule

module iob_dff(
	q,
	clk,
	rst,
	set_,
	en,
	d
	);
output	q;
input	clk;
input	rst,set_;
input	en;
input	d;
reg		q;
always @(posedge clk or posedge rst or negedge set_)
	if(~set_) q<=1;
	else if(rst) q<=0;
	else if(en) q<=d;
	else q<=q;
endmodule
/////////////////////////////////////////////////////////
//dff_n2mx & dff_2mx used in ILOGIC module
module dff_n2mx (
	q,
	clk,
	set_,
	rst,
	sel,
	sel_,
	init_b,
	in0,
	in1
	);
output	q;
input	clk,set_,rst;
input	sel,sel_,init_b;
input	in0,in1;

wire di =	({sel,sel_,init_b} == 3'b011) ? !in0 :
			({sel,sel_,init_b} == 3'b101) ? !in1 :
			({sel,sel_,init_b} == 3'b000) ? 1'b0 :
			({sel,sel_,init_b} == 3'b001) ? 1'b0 : 1'bx;
reg	qx;
always @(posedge clk or negedge set_ or posedge rst)
	if(~set_) qx <= 1;
	else if(rst) qx <= 0;
	else qx <= di;

assign q = ~qx;

endmodule

module dff_2mx (
	q,
	clk,
	set_,
	rst,
	sel,
	sel_,
	in0,
	in1
	);
output	q;
input	clk,set_,rst;
input	sel,sel_;
input	in0,in1;

wire di =	({sel,sel_} == 2'b01) ? !in0 :
			({sel,sel_} == 2'b10) ? !in1 : 1'bx;
reg	qx;
always @(posedge clk or negedge set_ or posedge rst)
	if(~set_) qx <= 1;
	else if(rst) qx <= 0;
	else qx <= di;

assign q = ~qx;

endmodule
//dff_2mx also used in OLOGIC module

//Updated 2015-06-09

//*************************************************
//Company:      CME
//Author:       hywang
//Filename:     fls_cbus.v
//Date:         20121225
//Function:     Serial flash controller control regiter
//*************************************************
`ifdef DLY
`else
`define DLY #1
`endif

module ahb_cfg_register (
                          clk, 
                          rst_n,
                          haddr,
                          htrans,
                          hwrite,
                          hwdata,
                          hrdata,
                          hready_out,
                          output_0,
                          output_1,
                          output_2,
                          output_3,
                          output_4,
                          output_5,
                          output_6,
                          output_7,
                          output_8,
                          output_9,
                          output_a
);      

parameter        ADDR0   =    8'h00,        
                 ADDR1   =    8'h04,        
                 ADDR2   =    8'h08,          
                 ADDR3   =    8'h0c,          
                 ADDR4   =    8'h10,        
                 ADDR5   =    8'h14, 
                 ADDR6   =    8'h18,
                 ADDR7   =    8'h1c,
                 ADDR8   =    8'h20,
                 ADDR9   =    8'h24,
                 ADDRA   =    8'h28;

//clock and reset
input          clk;
input          rst_n;

//PBUS slave/AS slave
input  [31:0]  haddr;
input  [1:0]   htrans;
input          hwrite;
input  [31:0]  hwdata;
output [31:0]  hrdata;
output         hready_out;
output [31:0]  output_0;
output [31:0]  output_1;
output [31:0]  output_2;
output [31:0]  output_3;
output [31:0]  output_4;
output [31:0]  output_5;
output [31:0]  output_6;
output [31:0]  output_7;
output [31:0]  output_8;
output [31:0]  output_9;
output [31:0]  output_a;

reg    [31:0]  hrdata;
reg    [31:0]  output_0;
reg    [31:0]  output_1;
reg    [31:0]  output_2;
reg    [31:0]  output_3;
reg    [31:0]  output_4;
reg    [31:0]  output_5;
reg    [31:0]  output_6;
reg    [31:0]  output_7;
reg    [31:0]  output_8;
reg    [31:0]  output_9;
reg    [31:0]  output_a;
//----------------------------------
wire   rd_req;
wire   wr_req;
reg    wr_en;
assign hready_out = 1;
assign rd_req = htrans[1] == 1 && hwrite == 0;
assign wr_req = htrans[1] == 1 && hwrite == 1;
always @(posedge clk or negedge rst_n) begin
    if(rst_n == 1'b0) begin
        wr_en        <= `DLY   1'h0;
    end
    else if(wr_req) begin
        wr_en        <= `DLY   1'h1;
    end
    else begin
        wr_en        <= `DLY   1'h0;
    end
end
always @(posedge clk or negedge rst_n) begin
    if(rst_n == 1'b0) begin
        hrdata        <= `DLY   1'h0;
    end
    else if(rd_req) begin
        case(haddr[7:0])  //n should be a necessary number 
            ADDR0 : hrdata        <= `DLY   output_0;
            ADDR1 : hrdata        <= `DLY   output_1;
            ADDR2 : hrdata        <= `DLY   output_2;
            ADDR3 : hrdata        <= `DLY   output_3;
            ADDR4 : hrdata        <= `DLY   output_4;
            ADDR5 : hrdata        <= `DLY   output_5;
            ADDR6 : hrdata        <= `DLY   output_6;
            ADDR7 : hrdata        <= `DLY   output_7;
            ADDR8 : hrdata        <= `DLY   output_8;
            ADDR9 : hrdata        <= `DLY   output_9;
            ADDRA : hrdata        <= `DLY   output_a;
          default : hrdata        <= `DLY   32'hdead_1234;
        endcase
    end
end
always @(posedge clk or negedge rst_n) begin
    if(rst_n == 1'b0) begin
        output_0        <= `DLY   32'h0;
        output_1        <= `DLY   32'h0;
        output_2        <= `DLY   32'h0;
        output_3        <= `DLY   32'h0;
        output_4        <= `DLY   32'h0;
        output_5        <= `DLY   32'h0;
        output_6        <= `DLY   32'h0;
        output_7        <= `DLY   32'h0;
        output_8        <= `DLY   32'h0;
        output_9        <= `DLY   32'h0;
        output_a        <= `DLY   32'h0;
    end
    else if(wr_en) begin
        case(haddr[7:0])  //n should be a necessary number 
            ADDR0 : output_0        <= `DLY   hwdata;
            ADDR1 : output_1        <= `DLY   hwdata;
            ADDR2 : output_2        <= `DLY   hwdata;
            ADDR3 : output_3        <= `DLY   hwdata;
            ADDR4 : output_4        <= `DLY   hwdata;
            ADDR5 : output_5        <= `DLY   hwdata;
            ADDR6 : output_6        <= `DLY   hwdata;
            ADDR7 : output_7        <= `DLY   hwdata;
            ADDR8 : output_8        <= `DLY   hwdata;
            ADDR9 : output_9        <= `DLY   hwdata;
            ADDRA : output_a        <= `DLY   hwdata;
          default : output_0        <= `DLY   output_0;
        endcase
    end
end



endmodule
       
// VPERL: GENERATED_BEG

module bus_top (
	cbi_pbus_addr,
	cbi_pbus_req,
	cbi_pbus_wdata,
	cbi_pbus_write,
	ctl_ahb_cfg_haddr_i,
	ctl_ahb_cfg_hburst_i,
	ctl_ahb_cfg_hready_i,
	ctl_ahb_cfg_hsel_i,
	ctl_ahb_cfg_hsize_i,
	ctl_ahb_cfg_htrans_i,
	ctl_ahb_cfg_hwdata_i,
	ctl_ahb_cfg_hwrite_i,
	hreg_haddr,
	hreg_htrans,
	hreg_hwdata,
	hreg_hwrite,
	o,
	pbus_gnt,
	pbus_rdata,
	pcsps_pbus_addr,
	pcsps_pbus_req,
	pcsps_pbus_wdata,
	pcsps_pbus_write,
	phy_ahb_haddr_i,
	phy_ahb_hburst_i,
	phy_ahb_hready_i,
	phy_ahb_hsel_i,
	phy_ahb_hsize_i,
	phy_ahb_htrans_i,
	phy_ahb_hwdata_i,
	phy_ahb_hwrite_i,
	cbi_pbus_gnt,
	cbi_pbus_rdata,
//	cfg_fp2ip_sel,
	clk_p,
	ctl_ahb_cfg_hrdata_o,
	ctl_ahb_cfg_hready_o,
	ctl_ahb_cfg_hresp_o,
	fp_cs_clk,
	fp_cs_rstn,
	hreg_hrdata,
	hreg_hready_out,
	i,
	pbus_addr,
	pbus_req,
	pbus_wdata,
	pbus_write,
	pclk_ddr,
	pcsps_pbus_gnt,
	pcsps_pbus_rdata,
	phy_ahb_hrdata_o,
	phy_ahb_hready_o,
	phy_ahb_hresp_o,
	s,
	usr_pbus_rstn 
);

output	[15:0]	cbi_pbus_addr;
output		cbi_pbus_req;
output	[31:0]	cbi_pbus_wdata;
output		cbi_pbus_write;
output	[31:0]	ctl_ahb_cfg_haddr_i;
output	[2:0]	ctl_ahb_cfg_hburst_i;
output		ctl_ahb_cfg_hready_i;
output		ctl_ahb_cfg_hsel_i;
output	[2:0]	ctl_ahb_cfg_hsize_i;
output	[1:0]	ctl_ahb_cfg_htrans_i;
output	[31:0]	ctl_ahb_cfg_hwdata_i;
output		ctl_ahb_cfg_hwrite_i;
output	[31:0]	hreg_haddr;
output	[1:0]	hreg_htrans;
output	[31:0]	hreg_hwdata;
output		hreg_hwrite;
output		o;
output		pbus_gnt;
output	[31:0]	pbus_rdata;
output	[15:0]	pcsps_pbus_addr;
output		pcsps_pbus_req;
output	[31:0]	pcsps_pbus_wdata;
output		pcsps_pbus_write;
output	[31:0]	phy_ahb_haddr_i;
output	[2:0]	phy_ahb_hburst_i;
output		phy_ahb_hready_i;
output		phy_ahb_hsel_i;
output	[2:0]	phy_ahb_hsize_i;
output	[1:0]	phy_ahb_htrans_i;
output	[31:0]	phy_ahb_hwdata_i;
output		phy_ahb_hwrite_i;
input		cbi_pbus_gnt;
input	[31:0]	cbi_pbus_rdata;
//input		cfg_fp2ip_sel;
input		clk_p;
input	[31:0]	ctl_ahb_cfg_hrdata_o;
input		ctl_ahb_cfg_hready_o;
input	[0:0]	ctl_ahb_cfg_hresp_o;
input		fp_cs_clk;
input		fp_cs_rstn;
input	[31:0]	hreg_hrdata;
input		hreg_hready_out;
input	[1:0]	i;
input	[31:0]	pbus_addr;
input		pbus_req;
input	[31:0]	pbus_wdata;
input		pbus_write;
input		pclk_ddr;
input		pcsps_pbus_gnt;
input	[31:0]	pcsps_pbus_rdata;
input	[31:0]	phy_ahb_hrdata_o;
input		phy_ahb_hready_o;
input	[0:0]	phy_ahb_hresp_o;
input		s;
input		usr_pbus_rstn;

parameter cfg_fp2ip_sel = 1'b0;

endmodule

// VPERL: GENERATED_END

module CFGMUX2S1_203 (
    i0,
    i1,
    o
`ifdef FM_HACK
	,SEL
`endif
);


input  [202:0] i0;
input  [202:0] i1;

output [202:0] o;

`ifdef CS_FORMALPRO_HACK
    wire          SEL;
`else
     `ifdef  SIMULATION
          reg  SEL = 1'b0;
     `else
		`ifdef FM_HACK
			input		SEL;
		`else
			parameter SEL = 1'b0;
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o =
                             SEL ? i1 :
                                   i0 ;
`endif
endmodule

module CFGMUX2S1_340 (
    i0,
    i1,
    o
`ifdef FM_HACK
	,SEL
`endif
);


input  [339:0] i0;
input  [339:0] i1;

output [339:0] o;

`ifdef CS_FORMALPRO_HACK
    wire          SEL;
`else
     `ifdef  SIMULATION
          reg  SEL = 1'b0;
     `else
		`ifdef FM_HACK
			input		SEL;
		`else
			parameter SEL = 1'b0;
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o =
                             SEL ? i1 :
                                   i0 ;
`endif
endmodule

module CFGMUX8S3_600 (
    i0,
    i1,
    i2,
    i3,
    i4,
    i5,
    i6,
    i7,
    o
`ifdef FM_HACK
	,SEL
`endif
);


input  [599:0] i0;
input  [599:0] i1;
input  [599:0] i2;
input  [599:0] i3;
input  [599:0] i4;
input  [599:0] i5;
input  [599:0] i6;
input  [599:0] i7;

output [599:0] o;

`ifdef CS_FORMALPRO_HACK
    wire [2:0]         SEL;
`else
     `ifdef  SIMULATION
          reg [2:0] SEL = 2'b00;
     `else
		`ifdef FM_HACK
			input	[2:0]	SEL;
		`else
			parameter SEL = 3'b000;
		`endif
     `endif
`endif

`ifndef CS_SW_SKEL
    assign         o =
                 (SEL == 3'b000) ? i0 :
                 (SEL == 3'b001) ? i1 :
                 (SEL == 3'b010) ? i2 :
                 (SEL == 3'b011) ? i3 :
                 (SEL == 3'b100) ? i4 :
                 (SEL == 3'b101) ? i5 :
                 (SEL == 3'b110) ? i6 :
                 (SEL == 3'b111) ? i7 : 1'bx;
`endif
endmodule

// VPERL: GENERATED_BEG

module ctrl_wrapper (
	ahb_cfg_hrdata_o,
	ahb_cfg_hready_o,
	ahb_cfg_hresp_o,
	dram_dfi_addr_p1,
	dram_dfi_addr_p0,
	dram_dfi_bank_p1,
	dram_dfi_bank_p0,
	dram_dfi_cas_n_p1,
	dram_dfi_cas_n_p0,
	dram_dfi_cke_p1,
	dram_dfi_cke_p0,
	dram_dfi_cs_n_duplicate_p1,
	dram_dfi_cs_n_duplicate_p0,
	dram_dfi_cs_n_p1,
	dram_dfi_cs_n_p0,
	dram_dfi_ctrlupd_req,
	dram_dfi_dram_clk_disable,
	dram_dfi_ecc_rddata_en_p1,
	dram_dfi_ecc_rddata_en_p0,
	dram_dfi_ecc_wrdata_en_p1,
	dram_dfi_ecc_wrdata_en_p0,
	dram_dfi_ecc_wrdata_p1,
	dram_dfi_ecc_wrdata_p0,
	dram_dfi_ecc_wrmask_p1,
	dram_dfi_ecc_wrmask_p0,
	dram_dfi_init_start,
	dram_dfi_ras_n_p1,
	dram_dfi_ras_n_p0,
	dram_dfi_rddata_en_p1,
	dram_dfi_rddata_en_p0,
	dram_dfi_rdlvl_delay,
	dram_dfi_rdlvl_delayn,
	dram_dfi_rdlvl_edge,
	dram_dfi_rdlvl_en,
	dram_dfi_rdlvl_gate_delay,
	dram_dfi_rdlvl_gate_en,
	dram_dfi_rdlvl_load,
	dram_dfi_reset_n_p1,
	dram_dfi_reset_n_p0,
	dram_dfi_we_n_p1,
	dram_dfi_we_n_p0,
	dram_dfi_wodt_p1,
	dram_dfi_wodt_p0,
	dram_dfi_wrdata_en_p1,
	dram_dfi_wrdata_en_p0,
	dram_dfi_wrdata_p1,
	dram_dfi_wrdata_p0,
	dram_dfi_wrlvl_delay,
	dram_dfi_wrlvl_en,
	dram_dfi_wrlvl_load,
	dram_dfi_wrlvl_strobe,
	dram_dfi_wrmask_p1,
	dram_dfi_wrmask_p0,
	gating_mc_clk,
	intr,
	o_p1,
	o_p0,
	r_ddr23phy_reg,
	r_system_pll_reg,
//	scan_ctl_o3,
//	scan_ctl_o2,
//	scan_ctl_o1,
//	scan_ctl_o0,
	ahb_cfg_haddr_i,
	ahb_cfg_hburst_i,
	ahb_cfg_hclk,
	ahb_cfg_hready_i,
	ahb_cfg_hresetn,
	ahb_cfg_hsel_i,
	ahb_cfg_hsize_i,
	ahb_cfg_htrans_i,
	ahb_cfg_hwdata_i,
	ahb_cfg_hwrite_i,
	axi_port02_aclk,
	axi_port02_arstn,
	axi_port00_aclk,
	axi_port00_arstn,
//	bus_ctl_sel,
	dram_dfi_ctrlupd_ack,
	dram_dfi_ecc_rddata_w1,
	dram_dfi_ecc_rddata_w0,
	dram_dfi_init_complete,
	dram_dfi_rddata_valid_w1,
	dram_dfi_rddata_valid_w0,
	dram_dfi_rddata_w1,
	dram_dfi_rddata_w0,
	dram_dfi_rdlvl_gate_mode,
	dram_dfi_rdlvl_mode,
	dram_dfi_rdlvl_resp,
	dram_dfi_wrlvl_mode,
	dram_dfi_wrlvl_resp,
	i_p1,
	i_p0,
	mc_clk,
	mc_rstn,
	ro_ddr23phy_reg
//	scan_ctl_i3,
//	scan_ctl_i2,
//	scan_ctl_i1,
//	scan_ctl_i0,
//	scan_en 
);

output	[31:0]	ahb_cfg_hrdata_o;
output		ahb_cfg_hready_o;
output	[1:0]	ahb_cfg_hresp_o;
output	[19:0]	dram_dfi_addr_p1;
output	[19:0]	dram_dfi_addr_p0;
output	[2:0]	dram_dfi_bank_p1;
output	[2:0]	dram_dfi_bank_p0;
output		dram_dfi_cas_n_p1;
output		dram_dfi_cas_n_p0;
output	[0:0]	dram_dfi_cke_p1;
output	[0:0]	dram_dfi_cke_p0;
output	[0:0]	dram_dfi_cs_n_duplicate_p1;
output	[0:0]	dram_dfi_cs_n_duplicate_p0;
output	[0:0]	dram_dfi_cs_n_p1;
output	[0:0]	dram_dfi_cs_n_p0;
output		dram_dfi_ctrlupd_req;
output		dram_dfi_dram_clk_disable;
output	[0:0]	dram_dfi_ecc_rddata_en_p1;
output	[0:0]	dram_dfi_ecc_rddata_en_p0;
output	[0:0]	dram_dfi_ecc_wrdata_en_p1;
output	[0:0]	dram_dfi_ecc_wrdata_en_p0;
output	[15:0]	dram_dfi_ecc_wrdata_p1;
output	[15:0]	dram_dfi_ecc_wrdata_p0;
output	[1:0]	dram_dfi_ecc_wrmask_p1;
output	[1:0]	dram_dfi_ecc_wrmask_p0;
output		dram_dfi_init_start;
output		dram_dfi_ras_n_p1;
output		dram_dfi_ras_n_p0;
output	[3:0]	dram_dfi_rddata_en_p1;
output	[3:0]	dram_dfi_rddata_en_p0;
output	[31:0]	dram_dfi_rdlvl_delay;
output	[31:0]	dram_dfi_rdlvl_delayn;
output	[0:0]	dram_dfi_rdlvl_edge;
output	[0:0]	dram_dfi_rdlvl_en;
output	[63:0]	dram_dfi_rdlvl_gate_delay;
output	[0:0]	dram_dfi_rdlvl_gate_en;
output	[0:0]	dram_dfi_rdlvl_load;
output		dram_dfi_reset_n_p1;
output		dram_dfi_reset_n_p0;
output		dram_dfi_we_n_p1;
output		dram_dfi_we_n_p0;
output	[0:0]	dram_dfi_wodt_p1;
output	[0:0]	dram_dfi_wodt_p0;
output	[3:0]	dram_dfi_wrdata_en_p1;
output	[3:0]	dram_dfi_wrdata_en_p0;
output	[63:0]	dram_dfi_wrdata_p1;
output	[63:0]	dram_dfi_wrdata_p0;
output	[31:0]	dram_dfi_wrlvl_delay;
output	[0:0]	dram_dfi_wrlvl_en;
output	[0:0]	dram_dfi_wrlvl_load;
output	[0:0]	dram_dfi_wrlvl_strobe;
output	[7:0]	dram_dfi_wrmask_p1;
output	[7:0]	dram_dfi_wrmask_p0;
output		gating_mc_clk;
output		intr;
output	[169:0]	o_p1;
output	[169:0]	o_p0;
output [2047:0]	r_ddr23phy_reg;
output	[31:0]	r_system_pll_reg;
input	[31:0]	ahb_cfg_haddr_i;
input	[2:0]	ahb_cfg_hburst_i;
input		ahb_cfg_hclk;
input		ahb_cfg_hready_i;
input		ahb_cfg_hresetn;
input		ahb_cfg_hsel_i;
input	[2:0]	ahb_cfg_hsize_i;
input	[1:0]	ahb_cfg_htrans_i;
input	[31:0]	ahb_cfg_hwdata_i;
input		ahb_cfg_hwrite_i;
input		axi_port02_aclk;
input		axi_port02_arstn;
input		axi_port00_aclk;
input		axi_port00_arstn;
//input		bus_ctl_sel;
input		dram_dfi_ctrlupd_ack;
input	[15:0]	dram_dfi_ecc_rddata_w1;
input	[15:0]	dram_dfi_ecc_rddata_w0;
input		dram_dfi_init_complete;
input	[3:0]	dram_dfi_rddata_valid_w1;
input	[3:0]	dram_dfi_rddata_valid_w0;
input	[63:0]	dram_dfi_rddata_w1;
input	[63:0]	dram_dfi_rddata_w0;
input	[1:0]	dram_dfi_rdlvl_gate_mode;
input	[1:0]	dram_dfi_rdlvl_mode;
input	[31:0]	dram_dfi_rdlvl_resp;
input	[1:0]	dram_dfi_wrlvl_mode;
input	[3:0]	dram_dfi_wrlvl_resp;
input	[279:0]	i_p1;
input	[279:0]	i_p0;
input		mc_clk;
input		mc_rstn;
input [2047:0]	ro_ddr23phy_reg;

parameter bus_ctl_sel = 1'b0;
parameter ddr_ctl_iso_en = 1'b0;
parameter ddr_ctl_pd = 1'b0;

endmodule

// VPERL: GENERATED_END

module DDR_CRG_CORE (
    x0_async_clk	,
    x1_async_clk	,
    mc_clk_us		,
    axi_port02_aclk     ,
    axi_port00_aclk     ,
    bypasspll_mc_clk_x4 ,
    mc_clk              ,
    pclk_ddr            ,
    axi_port02_arstn    ,
    axi_port00_arstn    ,
    mcfg_rstn           ,
    mc_rstn             ,
    rst_p_n             ,
    prstn_gx            ,
    fp_cs_clk           ,
    fp_cs_rstn          ,
    usr_pbus_rstn       ,
    pbus_rst_n          ,
    gating_mc_clk       ,
    r_system_pll_reg    ,
//    cfg_gx_soft_prst    ,
//    cfg_mc_bus_sel      ,
//    cfg_p0_sync         ,
//    cfg_p1_sync         ,
    p_rc                ,
    bypasspll_mc_clk_x4_ug,
    mc_clk_ug           ,
    axi_port00_aclk_ug  ,
    axi_port02_aclk_ug  ,
    axi_port00_aclk_us  ,
    axi_port02_aclk_us    
);
output		x0_async_clk	    ;
output		x1_async_clk	    ;	
output		mc_clk_us	    ;
output          axi_port02_aclk     ;
output          axi_port00_aclk     ;
output          bypasspll_mc_clk_x4 ;
output          mc_clk              ;
output          axi_port02_arstn    ;
output          axi_port00_arstn    ;
output          mcfg_rstn           ;//to reset ddr cfg reg only
output          mc_rstn             ;
input           fp_cs_clk           ;//clk to fp async bridge
output          fp_cs_rstn          ;//rst to fp async bridge
output          usr_pbus_rstn       ;//rst only reset the local pbus
output          rst_p_n             ;//rst from ccb to ddr
input           pclk_ddr            ;//pclk to the top reg
output          prstn_gx            ;//rst from ccb through ddr to gx
input           pbus_rst_n          ;

//input           cfg_gx_soft_prst    ;//from top.reg
input           gating_mc_clk       ; // default 0: ungate
//input           cfg_p0_sync         ;// 1: p0 sync to mc 0: async
//input           cfg_p1_sync         ;// 1: p1 sync to mc
//input           cfg_mc_bus_sel      ;
input   [31:0]  r_system_pll_reg    ;//ctrl bit from DDR own cfg domain; default 0

input           p_rc                ;
input           bypasspll_mc_clk_x4_ug;
input           mc_clk_ug           ;
input           axi_port00_aclk_ug  ;
input           axi_port02_aclk_ug  ;
input		axi_port00_aclk_us  ;
input  		axi_port02_aclk_us  ;

parameter cfg_gx_soft_prst = 1'b0;
parameter cfg_mc_bus_sel = 1'b0;


endmodule


module GX_CRG_CORE(
   // PCIE sii.cr
    pipe_clk,
    core_clk,
    core_clk_ug,
    aux_clk,
    aux_clk_g,
    pwr_rst_n,
    sticky_rst_n,
    non_sticky_rst_n,
    core_rst_n,
    pipe_rst_n,
    squelch_rst_n,
    aux_clk_active,

    resetB,
    clk_p,
    rst_p_n,
    pipe_glue_rstn,
    routing_pipe_glue_rstn,

    fp2HP_UsrRst_N,
    fp2HP_UsrRxRst_N,
    fp2HP_UsrTxRst_N,

    perst_n,
    pm_req_core_rst,
    pm_req_non_sticky_rst,
    pm_req_phy_rst,
    pm_req_sticky_rst,
    pm_sel_aux_clk,

    pclk_gx,//clk from ccb & through ddr
    prstn_gx,//rst from ccb & through ddr
    SERDES0_C0R0_CLK,

    mac_phy_rate,
    link_req_rst_not,
    SP2LP_pipe0_phystatus,
    fp_auxclk_sel_l12,
    cfg_pm_no_soft_rst,
    fp_pcie_only_rstn,
    app_ltssm_enable
);

input           pipe_clk;
output          core_clk;
output          core_clk_ug;

output          aux_clk;
output          aux_clk_g;
output          pwr_rst_n;
output          sticky_rst_n;
output          non_sticky_rst_n;
output          core_rst_n;
output          pipe_rst_n;
output          squelch_rst_n;
output          aux_clk_active;
output          resetB;
output          rst_p_n;
output          clk_p;
output          perst_n;
input           fp2HP_UsrRst_N;
input           fp2HP_UsrRxRst_N;
input           fp2HP_UsrTxRst_N;

input           pm_req_sticky_rst;
input           pm_req_core_rst;
input           pm_req_non_sticky_rst;
input           pm_sel_aux_clk;
input           pm_req_phy_rst;
input           routing_pipe_glue_rstn;
output          pipe_glue_rstn;

input           pclk_gx;//clk from ccb & through ddr
input           prstn_gx;//rst from ccb & through ddr

output  [0:0]   SERDES0_C0R0_CLK;

input           mac_phy_rate;
input           SP2LP_pipe0_phystatus;
input           link_req_rst_not;
input           fp_auxclk_sel_l12;
input           app_ltssm_enable;
input           cfg_pm_no_soft_rst;
input           fp_pcie_only_rstn;

parameter serdes_pd = 1'b0;

endmodule


module PCIE_V1 (
	SP2HP_L3RXClkCorUse,
	SP2HP_L3Rx8B10BDecMComDet,
	SP2HP_L3Rx8B10BDecPComDet,
	SP2HP_L3Rx8B10BUse,
	SP2HP_L3Rx8B10BUserDefCom,
	SP2HP_L3Rx8B10BValidComOnly,
	SP2HP_L3Rx4B5BAlignEn,
	SP2HP_L3Rx4B5BED,
	SP2HP_L3Rx4B5BSD,
	SP2HP_L3Rx4B5BUse,
	SP2HP_L3RxBitReverse,
	SP2HP_L3RxBufClr,
	SP2HP_L3RxBufDepth,
	SP2HP_L3RxBufUse,
	SP2HP_L3RxCAL10BEnable,
	SP2HP_L3RxCALAlignWord,
	SP2HP_L3RxCALDetUse,
	SP2HP_L3RxCALDouble,
	SP2HP_L3RxCALEnMComAlign,
	SP2HP_L3RxCALEnPComAlign,
	SP2HP_L3RxCALMComDet,
	SP2HP_L3RxCALMComValue,
	SP2HP_L3RxCALPComDet,
	SP2HP_L3RxCALPComValue,
	SP2HP_L3RxCALSlide,
	SP2HP_L3RxCALSlideMode,
	SP2HP_L3RxCHBondSeq1,
	SP2HP_L3RxCHBondSeq1En,
	SP2HP_L3RxCHBondSeq1Mask,
	SP2HP_L3RxClkCorAdjLen,
	SP2HP_L3RxClkCorSeq14,
	SP2HP_L3RxClkCorSeq13,
	SP2HP_L3RxClkCorSeq12,
	SP2HP_L3RxClkCorSeq11,
	SP2HP_L3RxClkCorSeq1En,
	SP2HP_L3RxDataWidth,
	SP2HP_L3RxGearboxADJSel,
	SP2HP_L3RxGearboxEnDec,
	SP2HP_L3RxGearboxSlip,
	SP2HP_L3RxGearboxUse,
	SP2HP_L3RxInternalWidth,
	SP2HP_L3RxLDEn,
	SP2HP_L3RxNELClkMuxSel,
	SP2HP_L3RxNLMux,
	SP2HP_L3RxNLMuxWidth,
	SP2HP_L3RxOOBBurstVal,
	SP2HP_L3RxOOBMaxBurst,
	SP2HP_L3RxOOBMaxCOMINIT,
	SP2HP_L3RxOOBMaxCOMSAS,
	SP2HP_L3RxOOBMaxCOMWAKE,
	SP2HP_L3RxOOBMinBurst,
	SP2HP_L3RxOOBMinCOMINIT,
	SP2HP_L3RxOOBMinCOMSAS,
	SP2HP_L3RxOOBMinCOMWAKE,
	SP2HP_L3RxOvrsmplEnAlign,
	SP2HP_L3RxOvrsmplMode,
	SP2HP_L3RxPMux,
	SP2HP_L3RxPRBSCntClr,
	SP2HP_L3RxPRBSTst,
	SP2HP_L3RxPRBSUsr,
	SP2HP_L3RxPRBSWidth,
	SP2HP_L3RxPRBSZCntClr,
	SP2HP_L3RxPolarity,
	SP2HP_L3RxRecClkMuxSel,
	SP2HP_L3RxSyncEn,
	SP2HP_L3RxSyncInvalidIncr,
	SP2HP_L3RxSyncThres,
	SP2HP_L3RxSyncThreshold,
	SP2HP_L3RxUClk2MuxSel,
	SP2HP_L3RxUClkMuxSel,
	SP2HP_L3Tx8B10BUse,
	SP2HP_L3Tx4B5BUse,
	SP2HP_L3TxBitReverse,
	SP2HP_L3TxBufClr,
	SP2HP_L3TxBufWidth,
	SP2HP_L3TxBufferUse,
	SP2HP_L3TxDMux,
	SP2HP_L3TxDataWidth,
	SP2HP_L3TxElecIdleAdj,
	SP2HP_L3TxFlMux,
	SP2HP_L3TxGearboxFunc,
	SP2HP_L3TxGearboxReadyPre,
	SP2HP_L3TxGearboxUse,
	SP2HP_L3TxInternalWidth,
	SP2HP_L3TxOOBMode,
	SP2HP_L3TxOutClkMuxSel,
	SP2HP_L3TxOvrsmplMode,
	SP2HP_L3TxPCIEBeaconPWidth,
	SP2HP_L3TxPCIEDetectRx,
	SP2HP_L3TxPCIEElecIdle,
	SP2HP_L3TxPClkMuxSel,
	SP2HP_L3TxPMux,
	SP2HP_L3TxPRBSErrCont,
	SP2HP_L3TxPRBSErrOne,
	SP2HP_L3TxPRBSTst,
	SP2HP_L3TxPRBSUsr,
	SP2HP_L3TxPRBSWidth,
	SP2HP_L3TxPolarity,
	SP2HP_L3TxSATAOOBComBurstVal,
	SP2HP_L3TxSATAOOBComRESET,
	SP2HP_L3TxSATAOOBComSAS,
	SP2HP_L3TxSATAOOBComWAKE,
	SP2HP_L3TxSATAOOBType,
	SP2HP_L3TxUClk2MuxSel,
	SP2HP_L3TxUClkMuxSel,
	SP2HP_L3TxUIASmpl,
	SP2HP_L3TxUsr8B10BDataK,
	SP2HP_L3TxUsr8B10BDispMode,
	SP2HP_L3TxUsr8B10BDispVal,
	SP2HP_L3TxUsrData,
	SP2HP_L3TxUsrGBHeader,
	SP2HP_L3TxUsrGBSequence,
	SP2HP_L3TxUsrGBStartSeq,
	SP2HP_L2RXClkCorUse,
	SP2HP_L2Rx8B10BDecMComDet,
	SP2HP_L2Rx8B10BDecPComDet,
	SP2HP_L2Rx8B10BUse,
	SP2HP_L2Rx8B10BUserDefCom,
	SP2HP_L2Rx8B10BValidComOnly,
	SP2HP_L2Rx4B5BAlignEn,
	SP2HP_L2Rx4B5BED,
	SP2HP_L2Rx4B5BSD,
	SP2HP_L2Rx4B5BUse,
	SP2HP_L2RxBitReverse,
	SP2HP_L2RxBufClr,
	SP2HP_L2RxBufDepth,
	SP2HP_L2RxBufUse,
	SP2HP_L2RxCAL10BEnable,
	SP2HP_L2RxCALAlignWord,
	SP2HP_L2RxCALDetUse,
	SP2HP_L2RxCALDouble,
	SP2HP_L2RxCALEnMComAlign,
	SP2HP_L2RxCALEnPComAlign,
	SP2HP_L2RxCALMComDet,
	SP2HP_L2RxCALMComValue,
	SP2HP_L2RxCALPComDet,
	SP2HP_L2RxCALPComValue,
	SP2HP_L2RxCALSlide,
	SP2HP_L2RxCALSlideMode,
	SP2HP_L2RxCHBondSeq1,
	SP2HP_L2RxCHBondSeq1En,
	SP2HP_L2RxCHBondSeq1Mask,
	SP2HP_L2RxClkCorAdjLen,
	SP2HP_L2RxClkCorSeq14,
	SP2HP_L2RxClkCorSeq13,
	SP2HP_L2RxClkCorSeq12,
	SP2HP_L2RxClkCorSeq11,
	SP2HP_L2RxClkCorSeq1En,
	SP2HP_L2RxDataWidth,
	SP2HP_L2RxGearboxADJSel,
	SP2HP_L2RxGearboxEnDec,
	SP2HP_L2RxGearboxSlip,
	SP2HP_L2RxGearboxUse,
	SP2HP_L2RxInternalWidth,
	SP2HP_L2RxLDEn,
	SP2HP_L2RxNELClkMuxSel,
	SP2HP_L2RxNLMux,
	SP2HP_L2RxNLMuxWidth,
	SP2HP_L2RxOOBBurstVal,
	SP2HP_L2RxOOBMaxBurst,
	SP2HP_L2RxOOBMaxCOMINIT,
	SP2HP_L2RxOOBMaxCOMSAS,
	SP2HP_L2RxOOBMaxCOMWAKE,
	SP2HP_L2RxOOBMinBurst,
	SP2HP_L2RxOOBMinCOMINIT,
	SP2HP_L2RxOOBMinCOMSAS,
	SP2HP_L2RxOOBMinCOMWAKE,
	SP2HP_L2RxOvrsmplEnAlign,
	SP2HP_L2RxOvrsmplMode,
	SP2HP_L2RxPMux,
	SP2HP_L2RxPRBSCntClr,
	SP2HP_L2RxPRBSTst,
	SP2HP_L2RxPRBSUsr,
	SP2HP_L2RxPRBSWidth,
	SP2HP_L2RxPRBSZCntClr,
	SP2HP_L2RxPolarity,
	SP2HP_L2RxRecClkMuxSel,
	SP2HP_L2RxSyncEn,
	SP2HP_L2RxSyncInvalidIncr,
	SP2HP_L2RxSyncThres,
	SP2HP_L2RxSyncThreshold,
	SP2HP_L2RxUClk2MuxSel,
	SP2HP_L2RxUClkMuxSel,
	SP2HP_L2Tx8B10BUse,
	SP2HP_L2Tx4B5BUse,
	SP2HP_L2TxBitReverse,
	SP2HP_L2TxBufClr,
	SP2HP_L2TxBufWidth,
	SP2HP_L2TxBufferUse,
	SP2HP_L2TxDMux,
	SP2HP_L2TxDataWidth,
	SP2HP_L2TxElecIdleAdj,
	SP2HP_L2TxFlMux,
	SP2HP_L2TxGearboxFunc,
	SP2HP_L2TxGearboxReadyPre,
	SP2HP_L2TxGearboxUse,
	SP2HP_L2TxInternalWidth,
	SP2HP_L2TxOOBMode,
	SP2HP_L2TxOutClkMuxSel,
	SP2HP_L2TxOvrsmplMode,
	SP2HP_L2TxPCIEBeaconPWidth,
	SP2HP_L2TxPCIEDetectRx,
	SP2HP_L2TxPCIEElecIdle,
	SP2HP_L2TxPClkMuxSel,
	SP2HP_L2TxPMux,
	SP2HP_L2TxPRBSErrCont,
	SP2HP_L2TxPRBSErrOne,
	SP2HP_L2TxPRBSTst,
	SP2HP_L2TxPRBSUsr,
	SP2HP_L2TxPRBSWidth,
	SP2HP_L2TxPolarity,
	SP2HP_L2TxSATAOOBComBurstVal,
	SP2HP_L2TxSATAOOBComRESET,
	SP2HP_L2TxSATAOOBComSAS,
	SP2HP_L2TxSATAOOBComWAKE,
	SP2HP_L2TxSATAOOBType,
	SP2HP_L2TxUClk2MuxSel,
	SP2HP_L2TxUClkMuxSel,
	SP2HP_L2TxUIASmpl,
	SP2HP_L2TxUsr8B10BDataK,
	SP2HP_L2TxUsr8B10BDispMode,
	SP2HP_L2TxUsr8B10BDispVal,
	SP2HP_L2TxUsrData,
	SP2HP_L2TxUsrGBHeader,
	SP2HP_L2TxUsrGBSequence,
	SP2HP_L2TxUsrGBStartSeq,
	SP2HP_L1RXClkCorUse,
	SP2HP_L1Rx8B10BDecMComDet,
	SP2HP_L1Rx8B10BDecPComDet,
	SP2HP_L1Rx8B10BUse,
	SP2HP_L1Rx8B10BUserDefCom,
	SP2HP_L1Rx8B10BValidComOnly,
	SP2HP_L1Rx4B5BAlignEn,
	SP2HP_L1Rx4B5BED,
	SP2HP_L1Rx4B5BSD,
	SP2HP_L1Rx4B5BUse,
	SP2HP_L1RxBitReverse,
	SP2HP_L1RxBufClr,
	SP2HP_L1RxBufDepth,
	SP2HP_L1RxBufUse,
	SP2HP_L1RxCAL10BEnable,
	SP2HP_L1RxCALAlignWord,
	SP2HP_L1RxCALDetUse,
	SP2HP_L1RxCALDouble,
	SP2HP_L1RxCALEnMComAlign,
	SP2HP_L1RxCALEnPComAlign,
	SP2HP_L1RxCALMComDet,
	SP2HP_L1RxCALMComValue,
	SP2HP_L1RxCALPComDet,
	SP2HP_L1RxCALPComValue,
	SP2HP_L1RxCALSlide,
	SP2HP_L1RxCALSlideMode,
	SP2HP_L1RxCHBondSeq1,
	SP2HP_L1RxCHBondSeq1En,
	SP2HP_L1RxCHBondSeq1Mask,
	SP2HP_L1RxClkCorAdjLen,
	SP2HP_L1RxClkCorSeq14,
	SP2HP_L1RxClkCorSeq13,
	SP2HP_L1RxClkCorSeq12,
	SP2HP_L1RxClkCorSeq11,
	SP2HP_L1RxClkCorSeq1En,
	SP2HP_L1RxDataWidth,
	SP2HP_L1RxGearboxADJSel,
	SP2HP_L1RxGearboxEnDec,
	SP2HP_L1RxGearboxSlip,
	SP2HP_L1RxGearboxUse,
	SP2HP_L1RxInternalWidth,
	SP2HP_L1RxLDEn,
	SP2HP_L1RxNELClkMuxSel,
	SP2HP_L1RxNLMux,
	SP2HP_L1RxNLMuxWidth,
	SP2HP_L1RxOOBBurstVal,
	SP2HP_L1RxOOBMaxBurst,
	SP2HP_L1RxOOBMaxCOMINIT,
	SP2HP_L1RxOOBMaxCOMSAS,
	SP2HP_L1RxOOBMaxCOMWAKE,
	SP2HP_L1RxOOBMinBurst,
	SP2HP_L1RxOOBMinCOMINIT,
	SP2HP_L1RxOOBMinCOMSAS,
	SP2HP_L1RxOOBMinCOMWAKE,
	SP2HP_L1RxOvrsmplEnAlign,
	SP2HP_L1RxOvrsmplMode,
	SP2HP_L1RxPMux,
	SP2HP_L1RxPRBSCntClr,
	SP2HP_L1RxPRBSTst,
	SP2HP_L1RxPRBSUsr,
	SP2HP_L1RxPRBSWidth,
	SP2HP_L1RxPRBSZCntClr,
	SP2HP_L1RxPolarity,
	SP2HP_L1RxRecClkMuxSel,
	SP2HP_L1RxSyncEn,
	SP2HP_L1RxSyncInvalidIncr,
	SP2HP_L1RxSyncThres,
	SP2HP_L1RxSyncThreshold,
	SP2HP_L1RxUClk2MuxSel,
	SP2HP_L1RxUClkMuxSel,
	SP2HP_L1Tx8B10BUse,
	SP2HP_L1Tx4B5BUse,
	SP2HP_L1TxBitReverse,
	SP2HP_L1TxBufClr,
	SP2HP_L1TxBufWidth,
	SP2HP_L1TxBufferUse,
	SP2HP_L1TxDMux,
	SP2HP_L1TxDataWidth,
	SP2HP_L1TxElecIdleAdj,
	SP2HP_L1TxFlMux,
	SP2HP_L1TxGearboxFunc,
	SP2HP_L1TxGearboxReadyPre,
	SP2HP_L1TxGearboxUse,
	SP2HP_L1TxInternalWidth,
	SP2HP_L1TxOOBMode,
	SP2HP_L1TxOutClkMuxSel,
	SP2HP_L1TxOvrsmplMode,
	SP2HP_L1TxPCIEBeaconPWidth,
	SP2HP_L1TxPCIEDetectRx,
	SP2HP_L1TxPCIEElecIdle,
	SP2HP_L1TxPClkMuxSel,
	SP2HP_L1TxPMux,
	SP2HP_L1TxPRBSErrCont,
	SP2HP_L1TxPRBSErrOne,
	SP2HP_L1TxPRBSTst,
	SP2HP_L1TxPRBSUsr,
	SP2HP_L1TxPRBSWidth,
	SP2HP_L1TxPolarity,
	SP2HP_L1TxSATAOOBComBurstVal,
	SP2HP_L1TxSATAOOBComRESET,
	SP2HP_L1TxSATAOOBComSAS,
	SP2HP_L1TxSATAOOBComWAKE,
	SP2HP_L1TxSATAOOBType,
	SP2HP_L1TxUClk2MuxSel,
	SP2HP_L1TxUClkMuxSel,
	SP2HP_L1TxUIASmpl,
	SP2HP_L1TxUsr8B10BDataK,
	SP2HP_L1TxUsr8B10BDispMode,
	SP2HP_L1TxUsr8B10BDispVal,
	SP2HP_L1TxUsrData,
	SP2HP_L1TxUsrGBHeader,
	SP2HP_L1TxUsrGBSequence,
	SP2HP_L1TxUsrGBStartSeq,
	SP2HP_L0RXClkCorUse,
	SP2HP_L0Rx8B10BDecMComDet,
	SP2HP_L0Rx8B10BDecPComDet,
	SP2HP_L0Rx8B10BUse,
	SP2HP_L0Rx8B10BUserDefCom,
	SP2HP_L0Rx8B10BValidComOnly,
	SP2HP_L0Rx4B5BAlignEn,
	SP2HP_L0Rx4B5BED,
	SP2HP_L0Rx4B5BSD,
	SP2HP_L0Rx4B5BUse,
	SP2HP_L0RxBitReverse,
	SP2HP_L0RxBufClr,
	SP2HP_L0RxBufDepth,
	SP2HP_L0RxBufUse,
	SP2HP_L0RxCAL10BEnable,
	SP2HP_L0RxCALAlignWord,
	SP2HP_L0RxCALDetUse,
	SP2HP_L0RxCALDouble,
	SP2HP_L0RxCALEnMComAlign,
	SP2HP_L0RxCALEnPComAlign,
	SP2HP_L0RxCALMComDet,
	SP2HP_L0RxCALMComValue,
	SP2HP_L0RxCALPComDet,
	SP2HP_L0RxCALPComValue,
	SP2HP_L0RxCALSlide,
	SP2HP_L0RxCALSlideMode,
	SP2HP_L0RxCHBondSeq1,
	SP2HP_L0RxCHBondSeq1En,
	SP2HP_L0RxCHBondSeq1Mask,
	SP2HP_L0RxClkCorAdjLen,
	SP2HP_L0RxClkCorSeq14,
	SP2HP_L0RxClkCorSeq13,
	SP2HP_L0RxClkCorSeq12,
	SP2HP_L0RxClkCorSeq11,
	SP2HP_L0RxClkCorSeq1En,
	SP2HP_L0RxDataWidth,
	SP2HP_L0RxGearboxADJSel,
	SP2HP_L0RxGearboxEnDec,
	SP2HP_L0RxGearboxSlip,
	SP2HP_L0RxGearboxUse,
	SP2HP_L0RxInternalWidth,
	SP2HP_L0RxLDEn,
	SP2HP_L0RxNELClkMuxSel,
	SP2HP_L0RxNLMux,
	SP2HP_L0RxNLMuxWidth,
	SP2HP_L0RxOOBBurstVal,
	SP2HP_L0RxOOBMaxBurst,
	SP2HP_L0RxOOBMaxCOMINIT,
	SP2HP_L0RxOOBMaxCOMSAS,
	SP2HP_L0RxOOBMaxCOMWAKE,
	SP2HP_L0RxOOBMinBurst,
	SP2HP_L0RxOOBMinCOMINIT,
	SP2HP_L0RxOOBMinCOMSAS,
	SP2HP_L0RxOOBMinCOMWAKE,
	SP2HP_L0RxOvrsmplEnAlign,
	SP2HP_L0RxOvrsmplMode,
	SP2HP_L0RxPMux,
	SP2HP_L0RxPRBSCntClr,
	SP2HP_L0RxPRBSTst,
	SP2HP_L0RxPRBSUsr,
	SP2HP_L0RxPRBSWidth,
	SP2HP_L0RxPRBSZCntClr,
	SP2HP_L0RxPolarity,
	SP2HP_L0RxRecClkMuxSel,
	SP2HP_L0RxSyncEn,
	SP2HP_L0RxSyncInvalidIncr,
	SP2HP_L0RxSyncThres,
	SP2HP_L0RxSyncThreshold,
	SP2HP_L0RxUClk2MuxSel,
	SP2HP_L0RxUClkMuxSel,
	SP2HP_L0Tx8B10BUse,
	SP2HP_L0Tx4B5BUse,
	SP2HP_L0TxBitReverse,
	SP2HP_L0TxBufClr,
	SP2HP_L0TxBufWidth,
	SP2HP_L0TxBufferUse,
	SP2HP_L0TxDMux,
	SP2HP_L0TxDataWidth,
	SP2HP_L0TxElecIdleAdj,
	SP2HP_L0TxFlMux,
	SP2HP_L0TxGearboxFunc,
	SP2HP_L0TxGearboxReadyPre,
	SP2HP_L0TxGearboxUse,
	SP2HP_L0TxInternalWidth,
	SP2HP_L0TxOOBMode,
	SP2HP_L0TxOutClkMuxSel,
	SP2HP_L0TxOvrsmplMode,
	SP2HP_L0TxPCIEBeaconPWidth,
	SP2HP_L0TxPCIEDetectRx,
	SP2HP_L0TxPCIEElecIdle,
	SP2HP_L0TxPClkMuxSel,
	SP2HP_L0TxPMux,
	SP2HP_L0TxPRBSErrCont,
	SP2HP_L0TxPRBSErrOne,
	SP2HP_L0TxPRBSTst,
	SP2HP_L0TxPRBSUsr,
	SP2HP_L0TxPRBSWidth,
	SP2HP_L0TxPolarity,
	SP2HP_L0TxSATAOOBComBurstVal,
	SP2HP_L0TxSATAOOBComRESET,
	SP2HP_L0TxSATAOOBComSAS,
	SP2HP_L0TxSATAOOBComWAKE,
	SP2HP_L0TxSATAOOBType,
	SP2HP_L0TxUClk2MuxSel,
	SP2HP_L0TxUClkMuxSel,
	SP2HP_L0TxUIASmpl,
	SP2HP_L0TxUsr8B10BDataK,
	SP2HP_L0TxUsr8B10BDispMode,
	SP2HP_L0TxUsr8B10BDispVal,
	SP2HP_L0TxUsrData,
	SP2HP_L0TxUsrGBHeader,
	SP2HP_L0TxUsrGBSequence,
	SP2HP_L0TxUsrGBStartSeq,
	SP2HP_LaneEn,
	SP2HP_PCIEMode,
	SP2HP_PonChgClkT2,
	SP2HP_PonChgClkT1,
	SP2HP_PonDfeCalT,
	SP2HP_PonInitT,
	SP2HP_PonOfstCalHiT,
	SP2HP_PonOfstCalLoT,
	SP2HP_PonPllDetT,
	SP2HP_PonPreDfeCalT,
	SP2HP_PonPrePllDetT,
	SP2HP_PonPreResCalT,
	SP2HP_PonPwrIntvalT,
	SP2HP_PonResCalHiT,
	SP2HP_PonResCalLoT,
	SP2HP_RxUnifClkSel,
	SP2HP_RxX4Mode,
	SP2HP_SSCEnX4,
	SP2HP_SysRstBSel,
	SP2HP_TxDetRxT4,
	SP2HP_TxDetRxT3,
	SP2HP_TxDetRxT2,
	SP2HP_TxDetRxT1,
	SP2HP_TxPhaseAlignT,
	SP2HP_TxX4Mode,
	SP2HP_UsrRst_N,
	SP2HP_UsrRxRst_N,
	SP2HP_UsrTxRst_N,
	SP2HP_xBG_SafeMode,
	SP2HP_xBG_pr200clkmux,
	SP2HP_xBG_pr100BRCal,
	SP2HP_xBG_pr100Rx,
	SP2HP_xBG_pr100Tx,
	SP2HP_xBG_pr100spare,
	SP2HP_xBG_prcal100Rx,
	SP2HP_xBG_prcal100Tx,
	SP2HP_xBG_prcal50Pll,
	SP2HP_xBG_prcal50spare,
	SP2HP_xBG_pwrdnB,
	SP2HP_xBG_trim,
	SP2HP_xCDR3_PIbiasTrim,
	SP2HP_xCDR3_PIcapTrim,
	SP2HP_xCDR3_PdivSelRx,
	SP2HP_xCDR3_SelFourFive,
	SP2HP_xCDR3_clkmode,
	SP2HP_xCDR3_dccen,
	SP2HP_xCDR3_dccfix,
	SP2HP_xCDR3_dcctrim,
	SP2HP_xCDR3_inc,
	SP2HP_xCDR3_incF,
	SP2HP_xCDR3_limHF,
	SP2HP_xCDR3_limLF,
	SP2HP_xCDR3_metamode,
	SP2HP_xCDR3_mult2F,
	SP2HP_xCDR3_offs,
	SP2HP_xCDR3_pwrdnB,
	SP2HP_xCDR3_updnsw,
	SP2HP_xCDR2_PIbiasTrim,
	SP2HP_xCDR2_PIcapTrim,
	SP2HP_xCDR2_PdivSelRx,
	SP2HP_xCDR2_SelFourFive,
	SP2HP_xCDR2_clkmode,
	SP2HP_xCDR2_dccen,
	SP2HP_xCDR2_dccfix,
	SP2HP_xCDR2_dcctrim,
	SP2HP_xCDR2_inc,
	SP2HP_xCDR2_incF,
	SP2HP_xCDR2_limHF,
	SP2HP_xCDR2_limLF,
	SP2HP_xCDR2_metamode,
	SP2HP_xCDR2_mult2F,
	SP2HP_xCDR2_offs,
	SP2HP_xCDR2_pwrdnB,
	SP2HP_xCDR2_updnsw,
	SP2HP_xCDR1_PIbiasTrim,
	SP2HP_xCDR1_PIcapTrim,
	SP2HP_xCDR1_PdivSelRx,
	SP2HP_xCDR1_SelFourFive,
	SP2HP_xCDR1_clkmode,
	SP2HP_xCDR1_dccen,
	SP2HP_xCDR1_dccfix,
	SP2HP_xCDR1_dcctrim,
	SP2HP_xCDR1_inc,
	SP2HP_xCDR1_incF,
	SP2HP_xCDR1_limHF,
	SP2HP_xCDR1_limLF,
	SP2HP_xCDR1_metamode,
	SP2HP_xCDR1_mult2F,
	SP2HP_xCDR1_offs,
	SP2HP_xCDR1_pwrdnB,
	SP2HP_xCDR1_updnsw,
	SP2HP_xCDR0_PIbiasTrim,
	SP2HP_xCDR0_PIcapTrim,
	SP2HP_xCDR0_PdivSelRx,
	SP2HP_xCDR0_SelFourFive,
	SP2HP_xCDR0_clkmode,
	SP2HP_xCDR0_dccen,
	SP2HP_xCDR0_dccfix,
	SP2HP_xCDR0_dcctrim,
	SP2HP_xCDR0_inc,
	SP2HP_xCDR0_incF,
	SP2HP_xCDR0_limHF,
	SP2HP_xCDR0_limLF,
	SP2HP_xCDR0_metamode,
	SP2HP_xCDR0_mult2F,
	SP2HP_xCDR0_offs,
	SP2HP_xCDR0_pwrdnB,
	SP2HP_xCDR0_updnsw,
	SP2HP_xCMU_clkmux_pwrdnB,
	SP2HP_xCMU_clkmux_swon,
	SP2HP_xCMU_cur_trim,
	SP2HP_xCMU_pwrdnB,
	SP2HP_xCMU_refclk_sel,
	SP2HP_xCTLE3_Adaps_En,
	SP2HP_xCTLE3_Adaps_inc,
	SP2HP_xCTLE3_memCap,
	SP2HP_xCTLE3_memRes3,
	SP2HP_xCTLE3_memRes2,
	SP2HP_xCTLE3_memRes1,
	SP2HP_xCTLE2_Adaps_En,
	SP2HP_xCTLE2_Adaps_inc,
	SP2HP_xCTLE2_memCap,
	SP2HP_xCTLE2_memRes3,
	SP2HP_xCTLE2_memRes2,
	SP2HP_xCTLE2_memRes1,
	SP2HP_xCTLE1_Adaps_En,
	SP2HP_xCTLE1_Adaps_inc,
	SP2HP_xCTLE1_memCap,
	SP2HP_xCTLE1_memRes3,
	SP2HP_xCTLE1_memRes2,
	SP2HP_xCTLE1_memRes1,
	SP2HP_xCTLE0_Adaps_En,
	SP2HP_xCTLE0_Adaps_inc,
	SP2HP_xCTLE0_memCap,
	SP2HP_xCTLE0_memRes3,
	SP2HP_xCTLE0_memRes2,
	SP2HP_xCTLE0_memRes1,
	SP2HP_xDFE3_Adaps_En,
	SP2HP_xDFE3_AnaClkEn,
	SP2HP_xDFE3_EyeScan_En,
	SP2HP_xDFE3_eqGain,
	SP2HP_xDFE3_isoGain,
	SP2HP_xDFE3_memDly,
	SP2HP_xDFE3_memTap4,
	SP2HP_xDFE3_memTap3,
	SP2HP_xDFE3_memTap2,
	SP2HP_xDFE3_memTap1,
	SP2HP_xDFE3_setDly,
	SP2HP_xDFE3_setEq,
	SP2HP_xDFE3_tapcursel,
	SP2HP_xDFE2_Adaps_En,
	SP2HP_xDFE2_AnaClkEn,
	SP2HP_xDFE2_EyeScan_En,
	SP2HP_xDFE2_eqGain,
	SP2HP_xDFE2_isoGain,
	SP2HP_xDFE2_memDly,
	SP2HP_xDFE2_memTap4,
	SP2HP_xDFE2_memTap3,
	SP2HP_xDFE2_memTap2,
	SP2HP_xDFE2_memTap1,
	SP2HP_xDFE2_setDly,
	SP2HP_xDFE2_setEq,
	SP2HP_xDFE2_tapcursel,
	SP2HP_xDFE1_Adaps_En,
	SP2HP_xDFE1_AnaClkEn,
	SP2HP_xDFE1_EyeScan_En,
	SP2HP_xDFE1_eqGain,
	SP2HP_xDFE1_isoGain,
	SP2HP_xDFE1_memDly,
	SP2HP_xDFE1_memTap4,
	SP2HP_xDFE1_memTap3,
	SP2HP_xDFE1_memTap2,
	SP2HP_xDFE1_memTap1,
	SP2HP_xDFE1_setDly,
	SP2HP_xDFE1_setEq,
	SP2HP_xDFE1_tapcursel,
	SP2HP_xDFE0_Adaps_En,
	SP2HP_xDFE0_AnaClkEn,
	SP2HP_xDFE0_EyeScan_En,
	SP2HP_xDFE0_eqGain,
	SP2HP_xDFE0_isoGain,
	SP2HP_xDFE0_memDly,
	SP2HP_xDFE0_memTap4,
	SP2HP_xDFE0_memTap3,
	SP2HP_xDFE0_memTap2,
	SP2HP_xDFE0_memTap1,
	SP2HP_xDFE0_setDly,
	SP2HP_xDFE0_setEq,
	SP2HP_xDFE0_tapcursel,
	SP2HP_xDFECalEn3_mem,
	SP2HP_xDFECalEn3_sel,
	SP2HP_xDFECalEn2_mem,
	SP2HP_xDFECalEn2_sel,
	SP2HP_xDFECalEn1_mem,
	SP2HP_xDFECalEn1_sel,
	SP2HP_xDFECalEn0_mem,
	SP2HP_xDFECalEn0_sel,
	SP2HP_xJTAG_AC_Signal,
	SP2HP_xJTAG_En,
	SP2HP_xJTAG_ShiftDR,
	SP2HP_xJTAG_acmode,
	SP2HP_xJTAG_ini_mem,
	SP2HP_xJTAG_pwrdnB,
	SP2HP_xJTAG_tap_resetB,
	SP2HP_xLane3_farlpbken,
	SP2HP_xLane3_nearlpbken,
	SP2HP_xLane2_farlpbken,
	SP2HP_xLane2_nearlpbken,
	SP2HP_xLane1_farlpbken,
	SP2HP_xLane1_nearlpbken,
	SP2HP_xLane0_farlpbken,
	SP2HP_xLane0_nearlpbken,
	SP2HP_xMisc_pwrdnB,
	SP2HP_xMisc_resetB,
	SP2HP_xOSC_CrntEn,
	SP2HP_xOSC_FSEn,
	SP2HP_xOSC_Rtrim,
	SP2HP_xOSC_pwrdnB,
	SP2HP_xOfstCal3_Ovrd,
	SP2HP_xOfstCal3_inc,
	SP2HP_xOfstCal3_mem,
	SP2HP_xOfstCal3_memCtrl,
	SP2HP_xOfstCal3_memEn,
	SP2HP_xOfstCal3_pwrdnB,
	SP2HP_xOfstCal2_Ovrd,
	SP2HP_xOfstCal2_inc,
	SP2HP_xOfstCal2_mem,
	SP2HP_xOfstCal2_memCtrl,
	SP2HP_xOfstCal2_memEn,
	SP2HP_xOfstCal2_pwrdnB,
	SP2HP_xOfstCal1_Ovrd,
	SP2HP_xOfstCal1_inc,
	SP2HP_xOfstCal1_mem,
	SP2HP_xOfstCal1_memCtrl,
	SP2HP_xOfstCal1_memEn,
	SP2HP_xOfstCal1_pwrdnB,
	SP2HP_xOfstCal0_Ovrd,
	SP2HP_xOfstCal0_inc,
	SP2HP_xOfstCal0_mem,
	SP2HP_xOfstCal0_memCtrl,
	SP2HP_xOfstCal0_memEn,
	SP2HP_xOfstCal0_pwrdnB,
	SP2HP_xPLL_CntlLimit_en,
	SP2HP_xPLL_FBDIV,
	SP2HP_xPLL_LockDet_Force_Lock,
	SP2HP_xPLL_Qpump_2,
	SP2HP_xPLL_Qpump_1,
	SP2HP_xPLL_REFDIV,
	SP2HP_xPLL_VCO_Ctuning,
	SP2HP_xPLL_buf_Itrim,
	SP2HP_xPLL_lockdet_en,
	SP2HP_xPLL_lockdet_period_sel,
	SP2HP_xPLL_lockdet_ppm_sel1,
	SP2HP_xPLL_lockdet_ppm_sel0,
	SP2HP_xPLL_pdivSel,
	SP2HP_xPLL_pwrdnB,
	SP2HP_xPLL_resetB,
	SP2HP_xPLL_selFourFive,
	SP2HP_xRX3_busdivSel,
	SP2HP_xRX3_pwrdnB,
	SP2HP_xRX3_set_phase,
	SP2HP_xRX3_slip_clk,
	SP2HP_xRX3_syncRxToUsrclk,
	SP2HP_xRX3_xrChicoOvrPh5to9,
	SP2HP_xRX3_xrChicoOvrd,
	SP2HP_xRX3_xrChicoOvrdEn,
	SP2HP_xRX2_busdivSel,
	SP2HP_xRX2_pwrdnB,
	SP2HP_xRX2_set_phase,
	SP2HP_xRX2_slip_clk,
	SP2HP_xRX2_syncRxToUsrclk,
	SP2HP_xRX2_xrChicoOvrPh5to9,
	SP2HP_xRX2_xrChicoOvrd,
	SP2HP_xRX2_xrChicoOvrdEn,
	SP2HP_xRX1_busdivSel,
	SP2HP_xRX1_pwrdnB,
	SP2HP_xRX1_set_phase,
	SP2HP_xRX1_slip_clk,
	SP2HP_xRX1_syncRxToUsrclk,
	SP2HP_xRX1_xrChicoOvrPh5to9,
	SP2HP_xRX1_xrChicoOvrd,
	SP2HP_xRX1_xrChicoOvrdEn,
	SP2HP_xRX0_busdivSel,
	SP2HP_xRX0_pwrdnB,
	SP2HP_xRX0_set_phase,
	SP2HP_xRX0_slip_clk,
	SP2HP_xRX0_syncRxToUsrclk,
	SP2HP_xRX0_xrChicoOvrPh5to9,
	SP2HP_xRX0_xrChicoOvrd,
	SP2HP_xRX0_xrChicoOvrdEn,
	SP2HP_xRXAFE3_InCMTrim,
	SP2HP_xRXAFE3_rcvShuntEn,
	SP2HP_xRXAFE3_rcvVssTermEn,
	SP2HP_xRXAFE3_rcvVttTermEn,
	SP2HP_xRXAFE3_termRes50En,
	SP2HP_xRXAFE2_InCMTrim,
	SP2HP_xRXAFE2_rcvShuntEn,
	SP2HP_xRXAFE2_rcvVssTermEn,
	SP2HP_xRXAFE2_rcvVttTermEn,
	SP2HP_xRXAFE2_termRes50En,
	SP2HP_xRXAFE1_InCMTrim,
	SP2HP_xRXAFE1_rcvShuntEn,
	SP2HP_xRXAFE1_rcvVssTermEn,
	SP2HP_xRXAFE1_rcvVttTermEn,
	SP2HP_xRXAFE1_termRes50En,
	SP2HP_xRXAFE0_InCMTrim,
	SP2HP_xRXAFE0_rcvShuntEn,
	SP2HP_xRXAFE0_rcvVssTermEn,
	SP2HP_xRXAFE0_rcvVttTermEn,
	SP2HP_xRXAFE0_termRes50En,
	SP2HP_xRXSquelch3_noSigLevel,
	SP2HP_xRXSquelch3_pwrdnB,
	SP2HP_xRXSquelch2_noSigLevel,
	SP2HP_xRXSquelch2_pwrdnB,
	SP2HP_xRXSquelch1_noSigLevel,
	SP2HP_xRXSquelch1_pwrdnB,
	SP2HP_xRXSquelch0_noSigLevel,
	SP2HP_xRXSquelch0_pwrdnB,
	SP2HP_xResCal_Bg_offset,
	SP2HP_xResCal_LPF_offset,
	SP2HP_xResCal_MemCtrl,
	SP2HP_xResCal_MemEn,
	SP2HP_xResCal_MemRes_Bg,
	SP2HP_xResCal_MemRes_LPF,
	SP2HP_xResCal_MemRes_Rx,
	SP2HP_xResCal_MemRes_Tx,
	SP2HP_xResCal_ResBg_sel,
	SP2HP_xResCal_ResLPF_sel,
	SP2HP_xResCal_ResRx_sel,
	SP2HP_xResCal_ResTx_sel,
	SP2HP_xResCal_Rx_offset,
	SP2HP_xResCal_Tx_offset,
	SP2HP_xTOP_DivOOB,
	SP2HP_xTOP_DivSSC,
	SP2HP_xTOP_DivSYS,
	SP2HP_xTOP_SYSClkSel,
	SP2HP_xTX3_ACCCLK_ROTATEH,
	SP2HP_xTX3_ACC_DIN_SEL,
	SP2HP_xTX3_ACC_NSEL,
	SP2HP_xTX3_ACC_OVERRIDE,
	SP2HP_xTX3_ACC_OVERRIDE_EN,
	SP2HP_xTX3_ACC_ROTATE,
	SP2HP_xTX3_ACC_UPDNSW,
	SP2HP_xTX3_Clk_pwrdnB,
	SP2HP_xTX3_DrvPostCursor,
	SP2HP_xTX3_DrvPreCursor,
	SP2HP_xTX3_Drv_pwrdnB,
	SP2HP_xTX3_Drvbiastrim,
	SP2HP_xTX3_Drvswing,
	SP2HP_xTX3_PI_captrim,
	SP2HP_xTX3_PI_pwrdnB,
	SP2HP_xTX3_PIbiasTrim,
	SP2HP_xTX3_Resl_En,
	SP2HP_xTX3_SSC_EN,
	SP2HP_xTX3_SSC_OVERRIDE,
	SP2HP_xTX3_SSC_OVERRIDE_EN,
	SP2HP_xTX3_SSC_TSEL,
	SP2HP_xTX3_Ser_pwrdnB,
	SP2HP_xTX3_Serbiastrim,
	SP2HP_xTX3_Vreftrim,
	SP2HP_xTX3_activepkEn,
	SP2HP_xTX3_busdivSel,
	SP2HP_xTX3_chico_cksel,
	SP2HP_xTX3_chico_pwrdnB,
	SP2HP_xTX3_ctune,
	SP2HP_xTX3_dccbiastrim,
	SP2HP_xTX3_dccerrtrim,
	SP2HP_xTX3_dccfix,
	SP2HP_xTX3_gmtune,
	SP2HP_xTX3_ovsdivEn,
	SP2HP_xTX3_pdivSel,
	SP2HP_xTX3_pwrdnB,
	SP2HP_xTX3_selFourFive,
	SP2HP_xTX3_sendidle,
	SP2HP_xTX3_syncTxToUsrclk,
	SP2HP_xTX3_tdccEn,
	SP2HP_xTX3_tdccovrd,
	SP2HP_xTX2_ACCCLK_ROTATEH,
	SP2HP_xTX2_ACC_DIN_SEL,
	SP2HP_xTX2_ACC_NSEL,
	SP2HP_xTX2_ACC_OVERRIDE,
	SP2HP_xTX2_ACC_OVERRIDE_EN,
	SP2HP_xTX2_ACC_ROTATE,
	SP2HP_xTX2_ACC_UPDNSW,
	SP2HP_xTX2_Clk_pwrdnB,
	SP2HP_xTX2_DrvPostCursor,
	SP2HP_xTX2_DrvPreCursor,
	SP2HP_xTX2_Drv_pwrdnB,
	SP2HP_xTX2_Drvbiastrim,
	SP2HP_xTX2_Drvswing,
	SP2HP_xTX2_PI_captrim,
	SP2HP_xTX2_PI_pwrdnB,
	SP2HP_xTX2_PIbiasTrim,
	SP2HP_xTX2_Resl_En,
	SP2HP_xTX2_SSC_EN,
	SP2HP_xTX2_SSC_OVERRIDE,
	SP2HP_xTX2_SSC_OVERRIDE_EN,
	SP2HP_xTX2_SSC_TSEL,
	SP2HP_xTX2_Ser_pwrdnB,
	SP2HP_xTX2_Serbiastrim,
	SP2HP_xTX2_Vreftrim,
	SP2HP_xTX2_activepkEn,
	SP2HP_xTX2_busdivSel,
	SP2HP_xTX2_chico_cksel,
	SP2HP_xTX2_chico_pwrdnB,
	SP2HP_xTX2_ctune,
	SP2HP_xTX2_dccbiastrim,
	SP2HP_xTX2_dccerrtrim,
	SP2HP_xTX2_dccfix,
	SP2HP_xTX2_gmtune,
	SP2HP_xTX2_ovsdivEn,
	SP2HP_xTX2_pdivSel,
	SP2HP_xTX2_pwrdnB,
	SP2HP_xTX2_selFourFive,
	SP2HP_xTX2_sendidle,
	SP2HP_xTX2_syncTxToUsrclk,
	SP2HP_xTX2_tdccEn,
	SP2HP_xTX2_tdccovrd,
	SP2HP_xTX1_ACCCLK_ROTATEH,
	SP2HP_xTX1_ACC_DIN_SEL,
	SP2HP_xTX1_ACC_NSEL,
	SP2HP_xTX1_ACC_OVERRIDE,
	SP2HP_xTX1_ACC_OVERRIDE_EN,
	SP2HP_xTX1_ACC_ROTATE,
	SP2HP_xTX1_ACC_UPDNSW,
	SP2HP_xTX1_Clk_pwrdnB,
	SP2HP_xTX1_DrvPostCursor,
	SP2HP_xTX1_DrvPreCursor,
	SP2HP_xTX1_Drv_pwrdnB,
	SP2HP_xTX1_Drvbiastrim,
	SP2HP_xTX1_Drvswing,
	SP2HP_xTX1_PI_captrim,
	SP2HP_xTX1_PI_pwrdnB,
	SP2HP_xTX1_PIbiasTrim,
	SP2HP_xTX1_Resl_En,
	SP2HP_xTX1_SSC_EN,
	SP2HP_xTX1_SSC_OVERRIDE,
	SP2HP_xTX1_SSC_OVERRIDE_EN,
	SP2HP_xTX1_SSC_TSEL,
	SP2HP_xTX1_Ser_pwrdnB,
	SP2HP_xTX1_Serbiastrim,
	SP2HP_xTX1_Vreftrim,
	SP2HP_xTX1_activepkEn,
	SP2HP_xTX1_busdivSel,
	SP2HP_xTX1_chico_cksel,
	SP2HP_xTX1_chico_pwrdnB,
	SP2HP_xTX1_ctune,
	SP2HP_xTX1_dccbiastrim,
	SP2HP_xTX1_dccerrtrim,
	SP2HP_xTX1_dccfix,
	SP2HP_xTX1_gmtune,
	SP2HP_xTX1_ovsdivEn,
	SP2HP_xTX1_pdivSel,
	SP2HP_xTX1_pwrdnB,
	SP2HP_xTX1_selFourFive,
	SP2HP_xTX1_sendidle,
	SP2HP_xTX1_syncTxToUsrclk,
	SP2HP_xTX1_tdccEn,
	SP2HP_xTX1_tdccovrd,
	SP2HP_xTX0_ACCCLK_ROTATEH,
	SP2HP_xTX0_ACC_DIN_SEL,
	SP2HP_xTX0_ACC_NSEL,
	SP2HP_xTX0_ACC_OVERRIDE,
	SP2HP_xTX0_ACC_OVERRIDE_EN,
	SP2HP_xTX0_ACC_ROTATE,
	SP2HP_xTX0_ACC_UPDNSW,
	SP2HP_xTX0_Clk_pwrdnB,
	SP2HP_xTX0_DrvPostCursor,
	SP2HP_xTX0_DrvPreCursor,
	SP2HP_xTX0_Drv_pwrdnB,
	SP2HP_xTX0_Drvbiastrim,
	SP2HP_xTX0_Drvswing,
	SP2HP_xTX0_PI_captrim,
	SP2HP_xTX0_PI_pwrdnB,
	SP2HP_xTX0_PIbiasTrim,
	SP2HP_xTX0_Resl_En,
	SP2HP_xTX0_SSC_EN,
	SP2HP_xTX0_SSC_OVERRIDE,
	SP2HP_xTX0_SSC_OVERRIDE_EN,
	SP2HP_xTX0_SSC_TSEL,
	SP2HP_xTX0_Ser_pwrdnB,
	SP2HP_xTX0_Serbiastrim,
	SP2HP_xTX0_Vreftrim,
	SP2HP_xTX0_activepkEn,
	SP2HP_xTX0_busdivSel,
	SP2HP_xTX0_chico_cksel,
	SP2HP_xTX0_chico_pwrdnB,
	SP2HP_xTX0_ctune,
	SP2HP_xTX0_dccbiastrim,
	SP2HP_xTX0_dccerrtrim,
	SP2HP_xTX0_dccfix,
	SP2HP_xTX0_gmtune,
	SP2HP_xTX0_ovsdivEn,
	SP2HP_xTX0_pdivSel,
	SP2HP_xTX0_pwrdnB,
	SP2HP_xTX0_selFourFive,
	SP2HP_xTX0_sendidle,
	SP2HP_xTX0_syncTxToUsrclk,
	SP2HP_xTX0_tdccEn,
	SP2HP_xTX0_tdccovrd,
	SP2HP_xTX_SSC_Align,
	SP2LP_pipe0_phystatus,
	app_parity_errs,
	aux_pm_en,
	cfg_2nd_reset,
	cfg_2ndbus_num,
	cfg_aer_int_msg_num,
	cfg_aer_rc_err_int,
	cfg_aer_rc_err_msi,
	cfg_atten_ind,
	cfg_bar5_limit,
	cfg_bar5_start,
	cfg_bar4_limit,
	cfg_bar4_start,
	cfg_bar3_limit,
	cfg_bar3_start,
	cfg_bar2_limit,
	cfg_bar2_start,
	cfg_bar1_limit,
	cfg_bar1_start,
	cfg_bar0_limit,
	cfg_bar0_start,
	cfg_bus_master_en,
	cfg_bw_mgt_int,
	cfg_eml_control,
	cfg_exp_rom_limit,
	cfg_exp_rom_start,
	cfg_int_disable,
	cfg_link_auto_bw_int,
	cfg_max_payload_size,
	cfg_max_rd_req_size,
	cfg_mem_space_en,
	cfg_msi_64,
	cfg_msi_addr,
	cfg_msi_data,
	cfg_msi_en,
	cfg_msi_mask,
	cfg_multi_msi_en,
	cfg_no_snoop_en,
	cfg_pbus_dev_num,
	cfg_pbus_num,
	cfg_pcie_cap_int_msg_num,
	cfg_pm_no_soft_rst,
	cfg_pme_int,
	cfg_pme_msi,
	cfg_pwr_ctrler_ctrl,
	cfg_pwr_ind,
	cfg_rcb,
	cfg_relax_order_en,
	cfg_send_cor_err,
	cfg_send_f_err,
	cfg_send_nf_err,
	cfg_subbus_num,
	cfg_sys_err_rc,
	clk_req_n,
	cxpl_debug_info,
	cxpl_debug_info_ei,
	diag_status_bus,
	en_aux_clk_g,
	hp_int,
	hp_msi,
	hp_pme,
	lbc_dbi_ack,
	lbc_dbi_dout,
	lbc_ext_addr,
	lbc_ext_bar_num,
	lbc_ext_cs,
	lbc_ext_dout,
	lbc_ext_io_access,
	lbc_ext_rom_access,
	lbc_ext_wr,
	link_req_rst_not,
	mac_phy_rate,
	mac_phy_rxstandby,
	pm_curnt_state,
	pm_dstate,
	pm_linkst_in_l2,
	pm_linkst_in_l1,
	pm_linkst_in_l0s,
	pm_linkst_l2_exit,
	pm_pme_en,
	pm_req_core_rst,
	pm_req_non_sticky_rst,
	pm_req_phy_rst,
	pm_req_sticky_rst,
	pm_sel_aux_clk,
	pm_status,
	pm_xtlh_block_tlp,
	radm_bypass_addr,
	radm_bypass_attr,
	radm_bypass_bcm,
	radm_bypass_byte_cnt,
	radm_bypass_cmpltr_id,
	radm_bypass_cpl_last,
	radm_bypass_cpl_status,
	radm_bypass_data,
	radm_bypass_dllp_abort,
	radm_bypass_dv,
	radm_bypass_dw_len,
	radm_bypass_dwen,
	radm_bypass_ecrc_err,
	radm_bypass_eot,
	radm_bypass_first_be,
	radm_bypass_fmt,
	radm_bypass_func_num,
	radm_bypass_hv,
	radm_bypass_in_membar_range,
	radm_bypass_io_req_in_range,
	radm_bypass_last_be,
	radm_bypass_poisoned,
	radm_bypass_reqid,
	radm_bypass_rom_in_range,
	radm_bypass_tag,
	radm_bypass_tc,
	radm_bypass_td,
	radm_bypass_tlp_abort,
	radm_bypass_type,
	radm_correctable_err,
	radm_cpl_timeout,
	radm_fatal_err,
	radm_grant_tlp_type,
	radm_inta_asserted,
	radm_inta_deasserted,
	radm_intb_asserted,
	radm_intb_deasserted,
	radm_intc_asserted,
	radm_intc_deasserted,
	radm_intd_asserted,
	radm_intd_deasserted,
	radm_msg_payload,
	radm_msg_req_id,
	radm_msg_unlock,
	radm_nonfatal_err,
	radm_pm_pme,
	radm_pm_to_ack,
	radm_pm_turnoff,
	radm_q_not_empty,
	radm_qoverflow,
	radm_timeout_cpl_attr,
	radm_timeout_cpl_len,
	radm_timeout_cpl_tag,
	radm_timeout_cpl_tc,
	radm_timeout_func_num,
	radm_trgt1_addr,
	radm_trgt1_attr,
	radm_trgt1_bcm,
	radm_trgt1_byte_cnt,
	radm_trgt1_cmpltr_id,
	radm_trgt1_cpl_last,
	radm_trgt1_cpl_status,
	radm_trgt1_data,
	radm_trgt1_dllp_abort,
	radm_trgt1_dv,
	radm_trgt1_dw_len,
	radm_trgt1_dwen,
	radm_trgt1_ecrc_err,
	radm_trgt1_eot,
	radm_trgt1_first_be,
	radm_trgt1_fmt,
	radm_trgt1_func_num,
	radm_trgt1_hv,
	radm_trgt1_in_membar_range,
	radm_trgt1_io_req_in_range,
	radm_trgt1_last_be,
	radm_trgt1_mem_type,
	radm_trgt1_poisoned,
	radm_trgt1_reqid,
	radm_trgt1_rom_in_range,
	radm_trgt1_tag,
	radm_trgt1_tc,
	radm_trgt1_td,
	radm_trgt1_tlp_abort,
	radm_trgt1_type,
	radm_vendor_msg,
	rdlh_link_up,
	routing_pipe_glue_rstn,
	rtlh_rfc_data,
	rtlh_rfc_upd,
	smlh_link_up,
	smlh_ltssm_state,
	smlh_req_rst_not,
	training_rst_n,
	trgt_cpl_timeout,
	trgt_lookup_empty,
	trgt_lookup_id,
	trgt_timeout_cpl_attr,
	trgt_timeout_cpl_func_num,
	trgt_timeout_cpl_len,
	trgt_timeout_cpl_tc,
	trgt_timeout_lookup_id,
	ven_msg_grant,
	ven_msi_grant,
	wake,
	xadm_client1_halt,
	xadm_client0_halt,
	xadm_cpld_cdts,
	xadm_cplh_cdts,
	xadm_npd_cdts,
	xadm_nph_cdts,
	xadm_pd_cdts,
	xadm_ph_cdts,
	HP2SP_L3RxCALDetected,
	HP2SP_L3RxGearboxIsSync,
	HP2SP_L3RxOOBCOMINITDet,
	HP2SP_L3RxOOBCOMSASDet,
	HP2SP_L3RxOOBCOMWAKEDet,
	HP2SP_L3RxOOBElecIdle,
	HP2SP_L3RxOvrsmplErr,
	HP2SP_L3RxPIPEPHYStatusRxDet,
	HP2SP_L3RxPIPERxDetected,
	HP2SP_L3RxPRBSErrCnt,
	HP2SP_L3RxPRBSZeroCnt,
	HP2SP_L3RxRecClk,
	HP2SP_L3RxRecClk2,
	HP2SP_L3RxSyncState,
	HP2SP_L3RxUsr8B10BDispErr,
	HP2SP_L3RxUsr8B10BEBCorCnt,
	HP2SP_L3RxUsr8B10BEBStat,
	HP2SP_L3RxUsr8B10BIsComma,
	HP2SP_L3RxUsr8B10BIsK,
	HP2SP_L3RxUsr8B10BNotInTable,
	HP2SP_L3RxUsr8B10BRunDisp,
	HP2SP_L3RxUsr8B10BValid,
	HP2SP_L3RxUsrData,
	HP2SP_L3RxUsrDataValid,
	HP2SP_L3RxUsrGBHeader,
	HP2SP_L3RxUsrGBHeaderValid,
	HP2SP_L3RxUsrGBStartSeq,
	HP2SP_L3TxBufStatus,
	HP2SP_L3TxOutClk,
	HP2SP_L3TxOutClk2,
	HP2SP_L3TxSATAOOBComFinish,
	HP2SP_L3TxUsrGBReady,
	HP2SP_L2RxCALDetected,
	HP2SP_L2RxGearboxIsSync,
	HP2SP_L2RxOOBCOMINITDet,
	HP2SP_L2RxOOBCOMSASDet,
	HP2SP_L2RxOOBCOMWAKEDet,
	HP2SP_L2RxOOBElecIdle,
	HP2SP_L2RxOvrsmplErr,
	HP2SP_L2RxPIPEPHYStatusRxDet,
	HP2SP_L2RxPIPERxDetected,
	HP2SP_L2RxPRBSErrCnt,
	HP2SP_L2RxPRBSZeroCnt,
	HP2SP_L2RxRecClk,
	HP2SP_L2RxRecClk2,
	HP2SP_L2RxSyncState,
	HP2SP_L2RxUsr8B10BDispErr,
	HP2SP_L2RxUsr8B10BEBCorCnt,
	HP2SP_L2RxUsr8B10BEBStat,
	HP2SP_L2RxUsr8B10BIsComma,
	HP2SP_L2RxUsr8B10BIsK,
	HP2SP_L2RxUsr8B10BNotInTable,
	HP2SP_L2RxUsr8B10BRunDisp,
	HP2SP_L2RxUsr8B10BValid,
	HP2SP_L2RxUsrData,
	HP2SP_L2RxUsrDataValid,
	HP2SP_L2RxUsrGBHeader,
	HP2SP_L2RxUsrGBHeaderValid,
	HP2SP_L2RxUsrGBStartSeq,
	HP2SP_L2TxBufStatus,
	HP2SP_L2TxOutClk,
	HP2SP_L2TxOutClk2,
	HP2SP_L2TxSATAOOBComFinish,
	HP2SP_L2TxUsrGBReady,
	HP2SP_L1RxCALDetected,
	HP2SP_L1RxGearboxIsSync,
	HP2SP_L1RxOOBCOMINITDet,
	HP2SP_L1RxOOBCOMSASDet,
	HP2SP_L1RxOOBCOMWAKEDet,
	HP2SP_L1RxOOBElecIdle,
	HP2SP_L1RxOvrsmplErr,
	HP2SP_L1RxPIPEPHYStatusRxDet,
	HP2SP_L1RxPIPERxDetected,
	HP2SP_L1RxPRBSErrCnt,
	HP2SP_L1RxPRBSZeroCnt,
	HP2SP_L1RxRecClk,
	HP2SP_L1RxRecClk2,
	HP2SP_L1RxSyncState,
	HP2SP_L1RxUsr8B10BDispErr,
	HP2SP_L1RxUsr8B10BEBCorCnt,
	HP2SP_L1RxUsr8B10BEBStat,
	HP2SP_L1RxUsr8B10BIsComma,
	HP2SP_L1RxUsr8B10BIsK,
	HP2SP_L1RxUsr8B10BNotInTable,
	HP2SP_L1RxUsr8B10BRunDisp,
	HP2SP_L1RxUsr8B10BValid,
	HP2SP_L1RxUsrData,
	HP2SP_L1RxUsrDataValid,
	HP2SP_L1RxUsrGBHeader,
	HP2SP_L1RxUsrGBHeaderValid,
	HP2SP_L1RxUsrGBStartSeq,
	HP2SP_L1TxBufStatus,
	HP2SP_L1TxOutClk,
	HP2SP_L1TxOutClk2,
	HP2SP_L1TxSATAOOBComFinish,
	HP2SP_L1TxUsrGBReady,
	HP2SP_L0RxCALDetected,
	HP2SP_L0RxGearboxIsSync,
	HP2SP_L0RxOOBCOMINITDet,
	HP2SP_L0RxOOBCOMSASDet,
	HP2SP_L0RxOOBCOMWAKEDet,
	HP2SP_L0RxOOBElecIdle,
	HP2SP_L0RxOvrsmplErr,
	HP2SP_L0RxPIPEPHYStatusRxDet,
	HP2SP_L0RxPIPERxDetected,
	HP2SP_L0RxPRBSErrCnt,
	HP2SP_L0RxPRBSZeroCnt,
	HP2SP_L0RxRecClk,
	HP2SP_L0RxRecClk2,
	HP2SP_L0RxSyncState,
	HP2SP_L0RxUsr8B10BDispErr,
	HP2SP_L0RxUsr8B10BEBCorCnt,
	HP2SP_L0RxUsr8B10BEBStat,
	HP2SP_L0RxUsr8B10BIsComma,
	HP2SP_L0RxUsr8B10BIsK,
	HP2SP_L0RxUsr8B10BNotInTable,
	HP2SP_L0RxUsr8B10BRunDisp,
	HP2SP_L0RxUsr8B10BValid,
	HP2SP_L0RxUsrData,
	HP2SP_L0RxUsrDataValid,
	HP2SP_L0RxUsrGBHeader,
	HP2SP_L0RxUsrGBHeaderValid,
	HP2SP_L0RxUsrGBStartSeq,
	HP2SP_L0TxBufStatus,
	HP2SP_L0TxOutClk,
	HP2SP_L0TxOutClk2,
	HP2SP_L0TxSATAOOBComFinish,
	HP2SP_L0TxUsrGBReady,
	HP2SP_PIPEPhyStatusForce,
	HP2SP_PIPEPhyStatusSoft,
	HP2SP_PowerOnDone,
	HP2SP_RxLDuAlignAcqr,
	HP2SP_SysClk,
	HP2SP_xPLL_DivClk,
	app_clk_req_n,
	app_cpld_ca,
	app_cplh_ca,
	app_err_advisory,
	app_err_bus,
	app_err_func_num,
	app_hdr_log,
	app_hdr_valid,
	app_init_rst,
	app_ltssm_enable,
	app_npd_ca,
	app_nph_ca,
	app_pd_ca,
	app_ph_ca,
	app_ready_entr_l23,
	app_req_entr_l1,
	app_req_exit_l1,
	app_req_retry_en,
	app_unlock_msg,
	app_xfer_pending,
	apps_pm_xmt_pme,
	apps_pm_xmt_turnoff,
	aux_clk,
	aux_clk_active,
	aux_clk_g,
	cfg_msi_pending,
	client1_addr_align_en,
	client1_cpl_bcm,
	client1_cpl_byte_cnt,
	client1_cpl_lookup_id,
	client1_cpl_status,
	client1_remote_req_id,
	client1_tlp_addr,
	client1_tlp_attr,
	client1_tlp_bad_eot,
	client1_tlp_byte_en,
	client1_tlp_byte_len,
	client1_tlp_data,
	client1_tlp_dv,
	client1_tlp_eot,
	client1_tlp_ep,
	client1_tlp_fmt,
	client1_tlp_func_num,
	client1_tlp_hv,
	client1_tlp_tc,
	client1_tlp_td,
	client1_tlp_tid,
	client1_tlp_type,
	client0_addr_align_en,
	client0_cpl_bcm,
	client0_cpl_byte_cnt,
	client0_cpl_lookup_id,
	client0_cpl_status,
	client0_remote_req_id,
	client0_tlp_addr,
	client0_tlp_attr,
	client0_tlp_bad_eot,
	client0_tlp_byte_en,
	client0_tlp_byte_len,
	client0_tlp_data,
	client0_tlp_dv,
	client0_tlp_eot,
	client0_tlp_ep,
	client0_tlp_fmt,
	client0_tlp_func_num,
	client0_tlp_hv,
	client0_tlp_tc,
	client0_tlp_td,
	client0_tlp_tid,
	client0_tlp_type,
	core_clk,
	core_clk_ug,
	core_rst_n,
	dbg_pba,
	dbg_table,
	fp_dbi_addr,
	fp_dbi_bar_num,
	fp_dbi_cs,
	fp_dbi_cs2,
	fp_dbi_din,
	fp_dbi_func_num,
	fp_dbi_io_access,
	fp_dbi_rom_access,
	fp_dbi_wr,
	ccb_dbi_addr,
	ccb_dbi_bar_num,
	ccb_dbi_cs,
	ccb_dbi_cs2,
	ccb_dbi_din,
	ccb_dbi_func_num,
	ccb_dbi_io_access,
	ccb_dbi_rom_access,
	ccb_dbi_wr,
	ccb_lbc_dbi_ack,
	ccb_lbc_dbi_dout,
	cbi_pbus_gnt,
	cbi_pbus_rdata,
	clk_p,
	rst_p_n,
	cbi_pbus_addr,
	cbi_pbus_write,
	cbi_pbus_req,
	cbi_pbus_wdata,
	device_type,
	diag_ctrl_bus,
	ext_lbc_ack,
	ext_lbc_din,
	fp2HP_pcs_usr_resetB,
	fp2LP_pipe_glue_rstn,
	non_sticky_rst_n,
	outband_pwrup_cmd,
	perst_n,
	phy_clk_req_n,
	pipe_clk,
	pipe_glue_rstn,
	pipe_rst_n,
	pwr_rst_n,
	rx_lane_flip_en,
	squelch_rst_n,
	sticky_rst_n,
	sys_atten_button_pressed,
	sys_aux_pwr_det,
	sys_cmd_cpled_int,
	sys_eml_interlock_engaged,
	sys_int,
	sys_mrl_sensor_chged,
	sys_mrl_sensor_state,
	sys_pre_det_chged,
	sys_pre_det_state,
	sys_pwr_fault_det,
	trgt1_radm_halt,
	trgt1_radm_pkt_halt,
	tx_lane_flip_en,
	ven_msg_attr,
	ven_msg_code,
	ven_msg_data,
	ven_msg_ep,
	ven_msg_fmt,
	ven_msg_func_num,
	ven_msg_len,
	ven_msg_req,
	ven_msg_tag,
	ven_msg_tc,
	ven_msg_td,
	ven_msg_type,
	ven_msi_func_num,
	ven_msi_req,
	ven_msi_tc,
	ven_msi_vector 
);

output		SP2HP_L3RXClkCorUse;
output		SP2HP_L3Rx8B10BDecMComDet;
output		SP2HP_L3Rx8B10BDecPComDet;
output		SP2HP_L3Rx8B10BUse;
output	[9:0]	SP2HP_L3Rx8B10BUserDefCom;
output		SP2HP_L3Rx8B10BValidComOnly;
output		SP2HP_L3Rx4B5BAlignEn;
output	[9:0]	SP2HP_L3Rx4B5BED;
output	[9:0]	SP2HP_L3Rx4B5BSD;
output		SP2HP_L3Rx4B5BUse;
output		SP2HP_L3RxBitReverse;
output		SP2HP_L3RxBufClr;
output	[1:0]	SP2HP_L3RxBufDepth;
output		SP2HP_L3RxBufUse;
output	[9:0]	SP2HP_L3RxCAL10BEnable;
output		SP2HP_L3RxCALAlignWord;
output		SP2HP_L3RxCALDetUse;
output		SP2HP_L3RxCALDouble;
output		SP2HP_L3RxCALEnMComAlign;
output		SP2HP_L3RxCALEnPComAlign;
output		SP2HP_L3RxCALMComDet;
output	[9:0]	SP2HP_L3RxCALMComValue;
output		SP2HP_L3RxCALPComDet;
output	[9:0]	SP2HP_L3RxCALPComValue;
output		SP2HP_L3RxCALSlide;
output	[1:0]	SP2HP_L3RxCALSlideMode;
output	[35:0]	SP2HP_L3RxCHBondSeq1;
output	[3:0]	SP2HP_L3RxCHBondSeq1En;
output	[8:0]	SP2HP_L3RxCHBondSeq1Mask;
output	[1:0]	SP2HP_L3RxClkCorAdjLen;
output	[8:0]	SP2HP_L3RxClkCorSeq14;
output	[8:0]	SP2HP_L3RxClkCorSeq13;
output	[8:0]	SP2HP_L3RxClkCorSeq12;
output	[8:0]	SP2HP_L3RxClkCorSeq11;
output	[3:0]	SP2HP_L3RxClkCorSeq1En;
output	[1:0]	SP2HP_L3RxDataWidth;
output		SP2HP_L3RxGearboxADJSel;
output		SP2HP_L3RxGearboxEnDec;
output		SP2HP_L3RxGearboxSlip;
output		SP2HP_L3RxGearboxUse;
output		SP2HP_L3RxInternalWidth;
output		SP2HP_L3RxLDEn;
output	[1:0]	SP2HP_L3RxNELClkMuxSel;
output	[1:0]	SP2HP_L3RxNLMux;
output		SP2HP_L3RxNLMuxWidth;
output	[2:0]	SP2HP_L3RxOOBBurstVal;
output	[5:0]	SP2HP_L3RxOOBMaxBurst;
output	[5:0]	SP2HP_L3RxOOBMaxCOMINIT;
output	[6:0]	SP2HP_L3RxOOBMaxCOMSAS;
output	[5:0]	SP2HP_L3RxOOBMaxCOMWAKE;
output	[5:0]	SP2HP_L3RxOOBMinBurst;
output	[5:0]	SP2HP_L3RxOOBMinCOMINIT;
output	[6:0]	SP2HP_L3RxOOBMinCOMSAS;
output	[5:0]	SP2HP_L3RxOOBMinCOMWAKE;
output		SP2HP_L3RxOvrsmplEnAlign;
output		SP2HP_L3RxOvrsmplMode;
output	[1:0]	SP2HP_L3RxPMux;
output		SP2HP_L3RxPRBSCntClr;
output	[2:0]	SP2HP_L3RxPRBSTst;
output	[39:0]	SP2HP_L3RxPRBSUsr;
output		SP2HP_L3RxPRBSWidth;
output		SP2HP_L3RxPRBSZCntClr;
output		SP2HP_L3RxPolarity;
output		SP2HP_L3RxRecClkMuxSel;
output		SP2HP_L3RxSyncEn;
output	[2:0]	SP2HP_L3RxSyncInvalidIncr;
output	[1:0]	SP2HP_L3RxSyncThres;
output	[2:0]	SP2HP_L3RxSyncThreshold;
output	[2:0]	SP2HP_L3RxUClk2MuxSel;
output	[1:0]	SP2HP_L3RxUClkMuxSel;
output		SP2HP_L3Tx8B10BUse;
output		SP2HP_L3Tx4B5BUse;
output		SP2HP_L3TxBitReverse;
output		SP2HP_L3TxBufClr;
output		SP2HP_L3TxBufWidth;
output		SP2HP_L3TxBufferUse;
output	[1:0]	SP2HP_L3TxDMux;
output	[1:0]	SP2HP_L3TxDataWidth;
output		SP2HP_L3TxElecIdleAdj;
output	[1:0]	SP2HP_L3TxFlMux;
output	[1:0]	SP2HP_L3TxGearboxFunc;
output	[2:0]	SP2HP_L3TxGearboxReadyPre;
output		SP2HP_L3TxGearboxUse;
output		SP2HP_L3TxInternalWidth;
output	[1:0]	SP2HP_L3TxOOBMode;
output	[1:0]	SP2HP_L3TxOutClkMuxSel;
output		SP2HP_L3TxOvrsmplMode;
output	[1:0]	SP2HP_L3TxPCIEBeaconPWidth;
output		SP2HP_L3TxPCIEDetectRx;
output		SP2HP_L3TxPCIEElecIdle;
output		SP2HP_L3TxPClkMuxSel;
output	[2:0]	SP2HP_L3TxPMux;
output		SP2HP_L3TxPRBSErrCont;
output		SP2HP_L3TxPRBSErrOne;
output	[2:0]	SP2HP_L3TxPRBSTst;
output	[39:0]	SP2HP_L3TxPRBSUsr;
output		SP2HP_L3TxPRBSWidth;
output		SP2HP_L3TxPolarity;
output	[3:0]	SP2HP_L3TxSATAOOBComBurstVal;
output		SP2HP_L3TxSATAOOBComRESET;
output		SP2HP_L3TxSATAOOBComSAS;
output		SP2HP_L3TxSATAOOBComWAKE;
output		SP2HP_L3TxSATAOOBType;
output	[1:0]	SP2HP_L3TxUClk2MuxSel;
output	[1:0]	SP2HP_L3TxUClkMuxSel;
output	[1:0]	SP2HP_L3TxUIASmpl;
output	[7:0]	SP2HP_L3TxUsr8B10BDataK;
output	[7:0]	SP2HP_L3TxUsr8B10BDispMode;
output	[7:0]	SP2HP_L3TxUsr8B10BDispVal;
output	[79:0]	SP2HP_L3TxUsrData;
output	[2:0]	SP2HP_L3TxUsrGBHeader;
output	[6:0]	SP2HP_L3TxUsrGBSequence;
output		SP2HP_L3TxUsrGBStartSeq;
output		SP2HP_L2RXClkCorUse;
output		SP2HP_L2Rx8B10BDecMComDet;
output		SP2HP_L2Rx8B10BDecPComDet;
output		SP2HP_L2Rx8B10BUse;
output	[9:0]	SP2HP_L2Rx8B10BUserDefCom;
output		SP2HP_L2Rx8B10BValidComOnly;
output		SP2HP_L2Rx4B5BAlignEn;
output	[9:0]	SP2HP_L2Rx4B5BED;
output	[9:0]	SP2HP_L2Rx4B5BSD;
output		SP2HP_L2Rx4B5BUse;
output		SP2HP_L2RxBitReverse;
output		SP2HP_L2RxBufClr;
output	[1:0]	SP2HP_L2RxBufDepth;
output		SP2HP_L2RxBufUse;
output	[9:0]	SP2HP_L2RxCAL10BEnable;
output		SP2HP_L2RxCALAlignWord;
output		SP2HP_L2RxCALDetUse;
output		SP2HP_L2RxCALDouble;
output		SP2HP_L2RxCALEnMComAlign;
output		SP2HP_L2RxCALEnPComAlign;
output		SP2HP_L2RxCALMComDet;
output	[9:0]	SP2HP_L2RxCALMComValue;
output		SP2HP_L2RxCALPComDet;
output	[9:0]	SP2HP_L2RxCALPComValue;
output		SP2HP_L2RxCALSlide;
output	[1:0]	SP2HP_L2RxCALSlideMode;
output	[35:0]	SP2HP_L2RxCHBondSeq1;
output	[3:0]	SP2HP_L2RxCHBondSeq1En;
output	[8:0]	SP2HP_L2RxCHBondSeq1Mask;
output	[1:0]	SP2HP_L2RxClkCorAdjLen;
output	[8:0]	SP2HP_L2RxClkCorSeq14;
output	[8:0]	SP2HP_L2RxClkCorSeq13;
output	[8:0]	SP2HP_L2RxClkCorSeq12;
output	[8:0]	SP2HP_L2RxClkCorSeq11;
output	[3:0]	SP2HP_L2RxClkCorSeq1En;
output	[1:0]	SP2HP_L2RxDataWidth;
output		SP2HP_L2RxGearboxADJSel;
output		SP2HP_L2RxGearboxEnDec;
output		SP2HP_L2RxGearboxSlip;
output		SP2HP_L2RxGearboxUse;
output		SP2HP_L2RxInternalWidth;
output		SP2HP_L2RxLDEn;
output	[1:0]	SP2HP_L2RxNELClkMuxSel;
output	[1:0]	SP2HP_L2RxNLMux;
output		SP2HP_L2RxNLMuxWidth;
output	[2:0]	SP2HP_L2RxOOBBurstVal;
output	[5:0]	SP2HP_L2RxOOBMaxBurst;
output	[5:0]	SP2HP_L2RxOOBMaxCOMINIT;
output	[6:0]	SP2HP_L2RxOOBMaxCOMSAS;
output	[5:0]	SP2HP_L2RxOOBMaxCOMWAKE;
output	[5:0]	SP2HP_L2RxOOBMinBurst;
output	[5:0]	SP2HP_L2RxOOBMinCOMINIT;
output	[6:0]	SP2HP_L2RxOOBMinCOMSAS;
output	[5:0]	SP2HP_L2RxOOBMinCOMWAKE;
output		SP2HP_L2RxOvrsmplEnAlign;
output		SP2HP_L2RxOvrsmplMode;
output	[1:0]	SP2HP_L2RxPMux;
output		SP2HP_L2RxPRBSCntClr;
output	[2:0]	SP2HP_L2RxPRBSTst;
output	[39:0]	SP2HP_L2RxPRBSUsr;
output		SP2HP_L2RxPRBSWidth;
output		SP2HP_L2RxPRBSZCntClr;
output		SP2HP_L2RxPolarity;
output		SP2HP_L2RxRecClkMuxSel;
output		SP2HP_L2RxSyncEn;
output	[2:0]	SP2HP_L2RxSyncInvalidIncr;
output	[1:0]	SP2HP_L2RxSyncThres;
output	[2:0]	SP2HP_L2RxSyncThreshold;
output	[2:0]	SP2HP_L2RxUClk2MuxSel;
output	[1:0]	SP2HP_L2RxUClkMuxSel;
output		SP2HP_L2Tx8B10BUse;
output		SP2HP_L2Tx4B5BUse;
output		SP2HP_L2TxBitReverse;
output		SP2HP_L2TxBufClr;
output		SP2HP_L2TxBufWidth;
output		SP2HP_L2TxBufferUse;
output	[1:0]	SP2HP_L2TxDMux;
output	[1:0]	SP2HP_L2TxDataWidth;
output		SP2HP_L2TxElecIdleAdj;
output	[1:0]	SP2HP_L2TxFlMux;
output	[1:0]	SP2HP_L2TxGearboxFunc;
output	[2:0]	SP2HP_L2TxGearboxReadyPre;
output		SP2HP_L2TxGearboxUse;
output		SP2HP_L2TxInternalWidth;
output	[1:0]	SP2HP_L2TxOOBMode;
output	[1:0]	SP2HP_L2TxOutClkMuxSel;
output		SP2HP_L2TxOvrsmplMode;
output	[1:0]	SP2HP_L2TxPCIEBeaconPWidth;
output		SP2HP_L2TxPCIEDetectRx;
output		SP2HP_L2TxPCIEElecIdle;
output		SP2HP_L2TxPClkMuxSel;
output	[2:0]	SP2HP_L2TxPMux;
output		SP2HP_L2TxPRBSErrCont;
output		SP2HP_L2TxPRBSErrOne;
output	[2:0]	SP2HP_L2TxPRBSTst;
output	[39:0]	SP2HP_L2TxPRBSUsr;
output		SP2HP_L2TxPRBSWidth;
output		SP2HP_L2TxPolarity;
output	[3:0]	SP2HP_L2TxSATAOOBComBurstVal;
output		SP2HP_L2TxSATAOOBComRESET;
output		SP2HP_L2TxSATAOOBComSAS;
output		SP2HP_L2TxSATAOOBComWAKE;
output		SP2HP_L2TxSATAOOBType;
output	[1:0]	SP2HP_L2TxUClk2MuxSel;
output	[1:0]	SP2HP_L2TxUClkMuxSel;
output	[1:0]	SP2HP_L2TxUIASmpl;
output	[7:0]	SP2HP_L2TxUsr8B10BDataK;
output	[7:0]	SP2HP_L2TxUsr8B10BDispMode;
output	[7:0]	SP2HP_L2TxUsr8B10BDispVal;
output	[79:0]	SP2HP_L2TxUsrData;
output	[2:0]	SP2HP_L2TxUsrGBHeader;
output	[6:0]	SP2HP_L2TxUsrGBSequence;
output		SP2HP_L2TxUsrGBStartSeq;
output		SP2HP_L1RXClkCorUse;
output		SP2HP_L1Rx8B10BDecMComDet;
output		SP2HP_L1Rx8B10BDecPComDet;
output		SP2HP_L1Rx8B10BUse;
output	[9:0]	SP2HP_L1Rx8B10BUserDefCom;
output		SP2HP_L1Rx8B10BValidComOnly;
output		SP2HP_L1Rx4B5BAlignEn;
output	[9:0]	SP2HP_L1Rx4B5BED;
output	[9:0]	SP2HP_L1Rx4B5BSD;
output		SP2HP_L1Rx4B5BUse;
output		SP2HP_L1RxBitReverse;
output		SP2HP_L1RxBufClr;
output	[1:0]	SP2HP_L1RxBufDepth;
output		SP2HP_L1RxBufUse;
output	[9:0]	SP2HP_L1RxCAL10BEnable;
output		SP2HP_L1RxCALAlignWord;
output		SP2HP_L1RxCALDetUse;
output		SP2HP_L1RxCALDouble;
output		SP2HP_L1RxCALEnMComAlign;
output		SP2HP_L1RxCALEnPComAlign;
output		SP2HP_L1RxCALMComDet;
output	[9:0]	SP2HP_L1RxCALMComValue;
output		SP2HP_L1RxCALPComDet;
output	[9:0]	SP2HP_L1RxCALPComValue;
output		SP2HP_L1RxCALSlide;
output	[1:0]	SP2HP_L1RxCALSlideMode;
output	[35:0]	SP2HP_L1RxCHBondSeq1;
output	[3:0]	SP2HP_L1RxCHBondSeq1En;
output	[8:0]	SP2HP_L1RxCHBondSeq1Mask;
output	[1:0]	SP2HP_L1RxClkCorAdjLen;
output	[8:0]	SP2HP_L1RxClkCorSeq14;
output	[8:0]	SP2HP_L1RxClkCorSeq13;
output	[8:0]	SP2HP_L1RxClkCorSeq12;
output	[8:0]	SP2HP_L1RxClkCorSeq11;
output	[3:0]	SP2HP_L1RxClkCorSeq1En;
output	[1:0]	SP2HP_L1RxDataWidth;
output		SP2HP_L1RxGearboxADJSel;
output		SP2HP_L1RxGearboxEnDec;
output		SP2HP_L1RxGearboxSlip;
output		SP2HP_L1RxGearboxUse;
output		SP2HP_L1RxInternalWidth;
output		SP2HP_L1RxLDEn;
output	[1:0]	SP2HP_L1RxNELClkMuxSel;
output	[1:0]	SP2HP_L1RxNLMux;
output		SP2HP_L1RxNLMuxWidth;
output	[2:0]	SP2HP_L1RxOOBBurstVal;
output	[5:0]	SP2HP_L1RxOOBMaxBurst;
output	[5:0]	SP2HP_L1RxOOBMaxCOMINIT;
output	[6:0]	SP2HP_L1RxOOBMaxCOMSAS;
output	[5:0]	SP2HP_L1RxOOBMaxCOMWAKE;
output	[5:0]	SP2HP_L1RxOOBMinBurst;
output	[5:0]	SP2HP_L1RxOOBMinCOMINIT;
output	[6:0]	SP2HP_L1RxOOBMinCOMSAS;
output	[5:0]	SP2HP_L1RxOOBMinCOMWAKE;
output		SP2HP_L1RxOvrsmplEnAlign;
output		SP2HP_L1RxOvrsmplMode;
output	[1:0]	SP2HP_L1RxPMux;
output		SP2HP_L1RxPRBSCntClr;
output	[2:0]	SP2HP_L1RxPRBSTst;
output	[39:0]	SP2HP_L1RxPRBSUsr;
output		SP2HP_L1RxPRBSWidth;
output		SP2HP_L1RxPRBSZCntClr;
output		SP2HP_L1RxPolarity;
output		SP2HP_L1RxRecClkMuxSel;
output		SP2HP_L1RxSyncEn;
output	[2:0]	SP2HP_L1RxSyncInvalidIncr;
output	[1:0]	SP2HP_L1RxSyncThres;
output	[2:0]	SP2HP_L1RxSyncThreshold;
output	[2:0]	SP2HP_L1RxUClk2MuxSel;
output	[1:0]	SP2HP_L1RxUClkMuxSel;
output		SP2HP_L1Tx8B10BUse;
output		SP2HP_L1Tx4B5BUse;
output		SP2HP_L1TxBitReverse;
output		SP2HP_L1TxBufClr;
output		SP2HP_L1TxBufWidth;
output		SP2HP_L1TxBufferUse;
output	[1:0]	SP2HP_L1TxDMux;
output	[1:0]	SP2HP_L1TxDataWidth;
output		SP2HP_L1TxElecIdleAdj;
output	[1:0]	SP2HP_L1TxFlMux;
output	[1:0]	SP2HP_L1TxGearboxFunc;
output	[2:0]	SP2HP_L1TxGearboxReadyPre;
output		SP2HP_L1TxGearboxUse;
output		SP2HP_L1TxInternalWidth;
output	[1:0]	SP2HP_L1TxOOBMode;
output	[1:0]	SP2HP_L1TxOutClkMuxSel;
output		SP2HP_L1TxOvrsmplMode;
output	[1:0]	SP2HP_L1TxPCIEBeaconPWidth;
output		SP2HP_L1TxPCIEDetectRx;
output		SP2HP_L1TxPCIEElecIdle;
output		SP2HP_L1TxPClkMuxSel;
output	[2:0]	SP2HP_L1TxPMux;
output		SP2HP_L1TxPRBSErrCont;
output		SP2HP_L1TxPRBSErrOne;
output	[2:0]	SP2HP_L1TxPRBSTst;
output	[39:0]	SP2HP_L1TxPRBSUsr;
output		SP2HP_L1TxPRBSWidth;
output		SP2HP_L1TxPolarity;
output	[3:0]	SP2HP_L1TxSATAOOBComBurstVal;
output		SP2HP_L1TxSATAOOBComRESET;
output		SP2HP_L1TxSATAOOBComSAS;
output		SP2HP_L1TxSATAOOBComWAKE;
output		SP2HP_L1TxSATAOOBType;
output	[1:0]	SP2HP_L1TxUClk2MuxSel;
output	[1:0]	SP2HP_L1TxUClkMuxSel;
output	[1:0]	SP2HP_L1TxUIASmpl;
output	[7:0]	SP2HP_L1TxUsr8B10BDataK;
output	[7:0]	SP2HP_L1TxUsr8B10BDispMode;
output	[7:0]	SP2HP_L1TxUsr8B10BDispVal;
output	[79:0]	SP2HP_L1TxUsrData;
output	[2:0]	SP2HP_L1TxUsrGBHeader;
output	[6:0]	SP2HP_L1TxUsrGBSequence;
output		SP2HP_L1TxUsrGBStartSeq;
output		SP2HP_L0RXClkCorUse;
output		SP2HP_L0Rx8B10BDecMComDet;
output		SP2HP_L0Rx8B10BDecPComDet;
output		SP2HP_L0Rx8B10BUse;
output	[9:0]	SP2HP_L0Rx8B10BUserDefCom;
output		SP2HP_L0Rx8B10BValidComOnly;
output		SP2HP_L0Rx4B5BAlignEn;
output	[9:0]	SP2HP_L0Rx4B5BED;
output	[9:0]	SP2HP_L0Rx4B5BSD;
output		SP2HP_L0Rx4B5BUse;
output		SP2HP_L0RxBitReverse;
output		SP2HP_L0RxBufClr;
output	[1:0]	SP2HP_L0RxBufDepth;
output		SP2HP_L0RxBufUse;
output	[9:0]	SP2HP_L0RxCAL10BEnable;
output		SP2HP_L0RxCALAlignWord;
output		SP2HP_L0RxCALDetUse;
output		SP2HP_L0RxCALDouble;
output		SP2HP_L0RxCALEnMComAlign;
output		SP2HP_L0RxCALEnPComAlign;
output		SP2HP_L0RxCALMComDet;
output	[9:0]	SP2HP_L0RxCALMComValue;
output		SP2HP_L0RxCALPComDet;
output	[9:0]	SP2HP_L0RxCALPComValue;
output		SP2HP_L0RxCALSlide;
output	[1:0]	SP2HP_L0RxCALSlideMode;
output	[35:0]	SP2HP_L0RxCHBondSeq1;
output	[3:0]	SP2HP_L0RxCHBondSeq1En;
output	[8:0]	SP2HP_L0RxCHBondSeq1Mask;
output	[1:0]	SP2HP_L0RxClkCorAdjLen;
output	[8:0]	SP2HP_L0RxClkCorSeq14;
output	[8:0]	SP2HP_L0RxClkCorSeq13;
output	[8:0]	SP2HP_L0RxClkCorSeq12;
output	[8:0]	SP2HP_L0RxClkCorSeq11;
output	[3:0]	SP2HP_L0RxClkCorSeq1En;
output	[1:0]	SP2HP_L0RxDataWidth;
output		SP2HP_L0RxGearboxADJSel;
output		SP2HP_L0RxGearboxEnDec;
output		SP2HP_L0RxGearboxSlip;
output		SP2HP_L0RxGearboxUse;
output		SP2HP_L0RxInternalWidth;
output		SP2HP_L0RxLDEn;
output	[1:0]	SP2HP_L0RxNELClkMuxSel;
output	[1:0]	SP2HP_L0RxNLMux;
output		SP2HP_L0RxNLMuxWidth;
output	[2:0]	SP2HP_L0RxOOBBurstVal;
output	[5:0]	SP2HP_L0RxOOBMaxBurst;
output	[5:0]	SP2HP_L0RxOOBMaxCOMINIT;
output	[6:0]	SP2HP_L0RxOOBMaxCOMSAS;
output	[5:0]	SP2HP_L0RxOOBMaxCOMWAKE;
output	[5:0]	SP2HP_L0RxOOBMinBurst;
output	[5:0]	SP2HP_L0RxOOBMinCOMINIT;
output	[6:0]	SP2HP_L0RxOOBMinCOMSAS;
output	[5:0]	SP2HP_L0RxOOBMinCOMWAKE;
output		SP2HP_L0RxOvrsmplEnAlign;
output		SP2HP_L0RxOvrsmplMode;
output	[1:0]	SP2HP_L0RxPMux;
output		SP2HP_L0RxPRBSCntClr;
output	[2:0]	SP2HP_L0RxPRBSTst;
output	[39:0]	SP2HP_L0RxPRBSUsr;
output		SP2HP_L0RxPRBSWidth;
output		SP2HP_L0RxPRBSZCntClr;
output		SP2HP_L0RxPolarity;
output		SP2HP_L0RxRecClkMuxSel;
output		SP2HP_L0RxSyncEn;
output	[2:0]	SP2HP_L0RxSyncInvalidIncr;
output	[1:0]	SP2HP_L0RxSyncThres;
output	[2:0]	SP2HP_L0RxSyncThreshold;
output	[2:0]	SP2HP_L0RxUClk2MuxSel;
output	[1:0]	SP2HP_L0RxUClkMuxSel;
output		SP2HP_L0Tx8B10BUse;
output		SP2HP_L0Tx4B5BUse;
output		SP2HP_L0TxBitReverse;
output		SP2HP_L0TxBufClr;
output		SP2HP_L0TxBufWidth;
output		SP2HP_L0TxBufferUse;
output	[1:0]	SP2HP_L0TxDMux;
output	[1:0]	SP2HP_L0TxDataWidth;
output		SP2HP_L0TxElecIdleAdj;
output	[1:0]	SP2HP_L0TxFlMux;
output	[1:0]	SP2HP_L0TxGearboxFunc;
output	[2:0]	SP2HP_L0TxGearboxReadyPre;
output		SP2HP_L0TxGearboxUse;
output		SP2HP_L0TxInternalWidth;
output	[1:0]	SP2HP_L0TxOOBMode;
output	[1:0]	SP2HP_L0TxOutClkMuxSel;
output		SP2HP_L0TxOvrsmplMode;
output	[1:0]	SP2HP_L0TxPCIEBeaconPWidth;
output		SP2HP_L0TxPCIEDetectRx;
output		SP2HP_L0TxPCIEElecIdle;
output		SP2HP_L0TxPClkMuxSel;
output	[2:0]	SP2HP_L0TxPMux;
output		SP2HP_L0TxPRBSErrCont;
output		SP2HP_L0TxPRBSErrOne;
output	[2:0]	SP2HP_L0TxPRBSTst;
output	[39:0]	SP2HP_L0TxPRBSUsr;
output		SP2HP_L0TxPRBSWidth;
output		SP2HP_L0TxPolarity;
output	[3:0]	SP2HP_L0TxSATAOOBComBurstVal;
output		SP2HP_L0TxSATAOOBComRESET;
output		SP2HP_L0TxSATAOOBComSAS;
output		SP2HP_L0TxSATAOOBComWAKE;
output		SP2HP_L0TxSATAOOBType;
output	[1:0]	SP2HP_L0TxUClk2MuxSel;
output	[1:0]	SP2HP_L0TxUClkMuxSel;
output	[1:0]	SP2HP_L0TxUIASmpl;
output	[7:0]	SP2HP_L0TxUsr8B10BDataK;
output	[7:0]	SP2HP_L0TxUsr8B10BDispMode;
output	[7:0]	SP2HP_L0TxUsr8B10BDispVal;
output	[79:0]	SP2HP_L0TxUsrData;
output	[2:0]	SP2HP_L0TxUsrGBHeader;
output	[6:0]	SP2HP_L0TxUsrGBSequence;
output		SP2HP_L0TxUsrGBStartSeq;
output	[3:0]	SP2HP_LaneEn;
output	[1:0]	SP2HP_PCIEMode;
output	[13:0]	SP2HP_PonChgClkT2;
output	[13:0]	SP2HP_PonChgClkT1;
output	[13:0]	SP2HP_PonDfeCalT;
output	[13:0]	SP2HP_PonInitT;
output	[13:0]	SP2HP_PonOfstCalHiT;
output	[13:0]	SP2HP_PonOfstCalLoT;
output	[13:0]	SP2HP_PonPllDetT;
output	[13:0]	SP2HP_PonPreDfeCalT;
output	[13:0]	SP2HP_PonPrePllDetT;
output	[13:0]	SP2HP_PonPreResCalT;
output	[13:0]	SP2HP_PonPwrIntvalT;
output	[13:0]	SP2HP_PonResCalHiT;
output	[13:0]	SP2HP_PonResCalLoT;
output	[3:0]	SP2HP_RxUnifClkSel;
output		SP2HP_RxX4Mode;
output		SP2HP_SSCEnX4;
output		SP2HP_SysRstBSel;
output	[6:0]	SP2HP_TxDetRxT4;
output	[2:0]	SP2HP_TxDetRxT3;
output	[2:0]	SP2HP_TxDetRxT2;
output	[5:0]	SP2HP_TxDetRxT1;
output	[13:0]	SP2HP_TxPhaseAlignT;
output		SP2HP_TxX4Mode;
output		SP2HP_UsrRst_N;
output		SP2HP_UsrRxRst_N;
output		SP2HP_UsrTxRst_N;
output		SP2HP_xBG_SafeMode;
output	[3:0]	SP2HP_xBG_pr200clkmux;
output	[3:0]	SP2HP_xBG_pr100BRCal;
output	[3:0]	SP2HP_xBG_pr100Rx;
output	[3:0]	SP2HP_xBG_pr100Tx;
output	[3:0]	SP2HP_xBG_pr100spare;
output	[3:0]	SP2HP_xBG_prcal100Rx;
output	[3:0]	SP2HP_xBG_prcal100Tx;
output	[1:0]	SP2HP_xBG_prcal50Pll;
output	[1:0]	SP2HP_xBG_prcal50spare;
output		SP2HP_xBG_pwrdnB;
output	[2:0]	SP2HP_xBG_trim;
output	[1:0]	SP2HP_xCDR3_PIbiasTrim;
output	[2:0]	SP2HP_xCDR3_PIcapTrim;
output	[1:0]	SP2HP_xCDR3_PdivSelRx;
output		SP2HP_xCDR3_SelFourFive;
output		SP2HP_xCDR3_clkmode;
output		SP2HP_xCDR3_dccen;
output		SP2HP_xCDR3_dccfix;
output		SP2HP_xCDR3_dcctrim;
output	[3:0]	SP2HP_xCDR3_inc;
output	[4:0]	SP2HP_xCDR3_incF;
output	[4:0]	SP2HP_xCDR3_limHF;
output	[4:0]	SP2HP_xCDR3_limLF;
output		SP2HP_xCDR3_metamode;
output		SP2HP_xCDR3_mult2F;
output	[7:0]	SP2HP_xCDR3_offs;
output		SP2HP_xCDR3_pwrdnB;
output		SP2HP_xCDR3_updnsw;
output	[1:0]	SP2HP_xCDR2_PIbiasTrim;
output	[2:0]	SP2HP_xCDR2_PIcapTrim;
output	[1:0]	SP2HP_xCDR2_PdivSelRx;
output		SP2HP_xCDR2_SelFourFive;
output		SP2HP_xCDR2_clkmode;
output		SP2HP_xCDR2_dccen;
output		SP2HP_xCDR2_dccfix;
output		SP2HP_xCDR2_dcctrim;
output	[3:0]	SP2HP_xCDR2_inc;
output	[4:0]	SP2HP_xCDR2_incF;
output	[4:0]	SP2HP_xCDR2_limHF;
output	[4:0]	SP2HP_xCDR2_limLF;
output		SP2HP_xCDR2_metamode;
output		SP2HP_xCDR2_mult2F;
output	[7:0]	SP2HP_xCDR2_offs;
output		SP2HP_xCDR2_pwrdnB;
output		SP2HP_xCDR2_updnsw;
output	[1:0]	SP2HP_xCDR1_PIbiasTrim;
output	[2:0]	SP2HP_xCDR1_PIcapTrim;
output	[1:0]	SP2HP_xCDR1_PdivSelRx;
output		SP2HP_xCDR1_SelFourFive;
output		SP2HP_xCDR1_clkmode;
output		SP2HP_xCDR1_dccen;
output		SP2HP_xCDR1_dccfix;
output		SP2HP_xCDR1_dcctrim;
output	[3:0]	SP2HP_xCDR1_inc;
output	[4:0]	SP2HP_xCDR1_incF;
output	[4:0]	SP2HP_xCDR1_limHF;
output	[4:0]	SP2HP_xCDR1_limLF;
output		SP2HP_xCDR1_metamode;
output		SP2HP_xCDR1_mult2F;
output	[7:0]	SP2HP_xCDR1_offs;
output		SP2HP_xCDR1_pwrdnB;
output		SP2HP_xCDR1_updnsw;
output	[1:0]	SP2HP_xCDR0_PIbiasTrim;
output	[2:0]	SP2HP_xCDR0_PIcapTrim;
output	[1:0]	SP2HP_xCDR0_PdivSelRx;
output		SP2HP_xCDR0_SelFourFive;
output		SP2HP_xCDR0_clkmode;
output		SP2HP_xCDR0_dccen;
output		SP2HP_xCDR0_dccfix;
output		SP2HP_xCDR0_dcctrim;
output	[3:0]	SP2HP_xCDR0_inc;
output	[4:0]	SP2HP_xCDR0_incF;
output	[4:0]	SP2HP_xCDR0_limHF;
output	[4:0]	SP2HP_xCDR0_limLF;
output		SP2HP_xCDR0_metamode;
output		SP2HP_xCDR0_mult2F;
output	[7:0]	SP2HP_xCDR0_offs;
output		SP2HP_xCDR0_pwrdnB;
output		SP2HP_xCDR0_updnsw;
output		SP2HP_xCMU_clkmux_pwrdnB;
output		SP2HP_xCMU_clkmux_swon;
output	[1:0]	SP2HP_xCMU_cur_trim;
output		SP2HP_xCMU_pwrdnB;
output	[5:0]	SP2HP_xCMU_refclk_sel;
output		SP2HP_xCTLE3_Adaps_En;
output	[1:0]	SP2HP_xCTLE3_Adaps_inc;
output	[3:0]	SP2HP_xCTLE3_memCap;
output	[2:0]	SP2HP_xCTLE3_memRes3;
output	[1:0]	SP2HP_xCTLE3_memRes2;
output	[1:0]	SP2HP_xCTLE3_memRes1;
output		SP2HP_xCTLE2_Adaps_En;
output	[1:0]	SP2HP_xCTLE2_Adaps_inc;
output	[3:0]	SP2HP_xCTLE2_memCap;
output	[2:0]	SP2HP_xCTLE2_memRes3;
output	[1:0]	SP2HP_xCTLE2_memRes2;
output	[1:0]	SP2HP_xCTLE2_memRes1;
output		SP2HP_xCTLE1_Adaps_En;
output	[1:0]	SP2HP_xCTLE1_Adaps_inc;
output	[3:0]	SP2HP_xCTLE1_memCap;
output	[2:0]	SP2HP_xCTLE1_memRes3;
output	[1:0]	SP2HP_xCTLE1_memRes2;
output	[1:0]	SP2HP_xCTLE1_memRes1;
output		SP2HP_xCTLE0_Adaps_En;
output	[1:0]	SP2HP_xCTLE0_Adaps_inc;
output	[3:0]	SP2HP_xCTLE0_memCap;
output	[2:0]	SP2HP_xCTLE0_memRes3;
output	[1:0]	SP2HP_xCTLE0_memRes2;
output	[1:0]	SP2HP_xCTLE0_memRes1;
output		SP2HP_xDFE3_Adaps_En;
output		SP2HP_xDFE3_AnaClkEn;
output		SP2HP_xDFE3_EyeScan_En;
output	[4:0]	SP2HP_xDFE3_eqGain;
output	[2:0]	SP2HP_xDFE3_isoGain;
output	[5:0]	SP2HP_xDFE3_memDly;
output	[3:0]	SP2HP_xDFE3_memTap4;
output	[3:0]	SP2HP_xDFE3_memTap3;
output	[4:0]	SP2HP_xDFE3_memTap2;
output	[4:0]	SP2HP_xDFE3_memTap1;
output		SP2HP_xDFE3_setDly;
output		SP2HP_xDFE3_setEq;
output		SP2HP_xDFE3_tapcursel;
output		SP2HP_xDFE2_Adaps_En;
output		SP2HP_xDFE2_AnaClkEn;
output		SP2HP_xDFE2_EyeScan_En;
output	[4:0]	SP2HP_xDFE2_eqGain;
output	[2:0]	SP2HP_xDFE2_isoGain;
output	[5:0]	SP2HP_xDFE2_memDly;
output	[3:0]	SP2HP_xDFE2_memTap4;
output	[3:0]	SP2HP_xDFE2_memTap3;
output	[4:0]	SP2HP_xDFE2_memTap2;
output	[4:0]	SP2HP_xDFE2_memTap1;
output		SP2HP_xDFE2_setDly;
output		SP2HP_xDFE2_setEq;
output		SP2HP_xDFE2_tapcursel;
output		SP2HP_xDFE1_Adaps_En;
output		SP2HP_xDFE1_AnaClkEn;
output		SP2HP_xDFE1_EyeScan_En;
output	[4:0]	SP2HP_xDFE1_eqGain;
output	[2:0]	SP2HP_xDFE1_isoGain;
output	[5:0]	SP2HP_xDFE1_memDly;
output	[3:0]	SP2HP_xDFE1_memTap4;
output	[3:0]	SP2HP_xDFE1_memTap3;
output	[4:0]	SP2HP_xDFE1_memTap2;
output	[4:0]	SP2HP_xDFE1_memTap1;
output		SP2HP_xDFE1_setDly;
output		SP2HP_xDFE1_setEq;
output		SP2HP_xDFE1_tapcursel;
output		SP2HP_xDFE0_Adaps_En;
output		SP2HP_xDFE0_AnaClkEn;
output		SP2HP_xDFE0_EyeScan_En;
output	[4:0]	SP2HP_xDFE0_eqGain;
output	[2:0]	SP2HP_xDFE0_isoGain;
output	[5:0]	SP2HP_xDFE0_memDly;
output	[3:0]	SP2HP_xDFE0_memTap4;
output	[3:0]	SP2HP_xDFE0_memTap3;
output	[4:0]	SP2HP_xDFE0_memTap2;
output	[4:0]	SP2HP_xDFE0_memTap1;
output		SP2HP_xDFE0_setDly;
output		SP2HP_xDFE0_setEq;
output		SP2HP_xDFE0_tapcursel;
output		SP2HP_xDFECalEn3_mem;
output		SP2HP_xDFECalEn3_sel;
output		SP2HP_xDFECalEn2_mem;
output		SP2HP_xDFECalEn2_sel;
output		SP2HP_xDFECalEn1_mem;
output		SP2HP_xDFECalEn1_sel;
output		SP2HP_xDFECalEn0_mem;
output		SP2HP_xDFECalEn0_sel;
output		SP2HP_xJTAG_AC_Signal;
output		SP2HP_xJTAG_En;
output		SP2HP_xJTAG_ShiftDR;
output		SP2HP_xJTAG_acmode;
output		SP2HP_xJTAG_ini_mem;
output		SP2HP_xJTAG_pwrdnB;
output		SP2HP_xJTAG_tap_resetB;
output		SP2HP_xLane3_farlpbken;
output		SP2HP_xLane3_nearlpbken;
output		SP2HP_xLane2_farlpbken;
output		SP2HP_xLane2_nearlpbken;
output		SP2HP_xLane1_farlpbken;
output		SP2HP_xLane1_nearlpbken;
output		SP2HP_xLane0_farlpbken;
output		SP2HP_xLane0_nearlpbken;
output		SP2HP_xMisc_pwrdnB;
output		SP2HP_xMisc_resetB;
output		SP2HP_xOSC_CrntEn;
output		SP2HP_xOSC_FSEn;
output	[3:0]	SP2HP_xOSC_Rtrim;
output		SP2HP_xOSC_pwrdnB;
output		SP2HP_xOfstCal3_Ovrd;
output	[1:0]	SP2HP_xOfstCal3_inc;
output	[4:0]	SP2HP_xOfstCal3_mem;
output		SP2HP_xOfstCal3_memCtrl;
output		SP2HP_xOfstCal3_memEn;
output		SP2HP_xOfstCal3_pwrdnB;
output		SP2HP_xOfstCal2_Ovrd;
output	[1:0]	SP2HP_xOfstCal2_inc;
output	[4:0]	SP2HP_xOfstCal2_mem;
output		SP2HP_xOfstCal2_memCtrl;
output		SP2HP_xOfstCal2_memEn;
output		SP2HP_xOfstCal2_pwrdnB;
output		SP2HP_xOfstCal1_Ovrd;
output	[1:0]	SP2HP_xOfstCal1_inc;
output	[4:0]	SP2HP_xOfstCal1_mem;
output		SP2HP_xOfstCal1_memCtrl;
output		SP2HP_xOfstCal1_memEn;
output		SP2HP_xOfstCal1_pwrdnB;
output		SP2HP_xOfstCal0_Ovrd;
output	[1:0]	SP2HP_xOfstCal0_inc;
output	[4:0]	SP2HP_xOfstCal0_mem;
output		SP2HP_xOfstCal0_memCtrl;
output		SP2HP_xOfstCal0_memEn;
output		SP2HP_xOfstCal0_pwrdnB;
output		SP2HP_xPLL_CntlLimit_en;
output	[5:0]	SP2HP_xPLL_FBDIV;
output		SP2HP_xPLL_LockDet_Force_Lock;
output	[3:0]	SP2HP_xPLL_Qpump_2;
output	[3:0]	SP2HP_xPLL_Qpump_1;
output	[5:0]	SP2HP_xPLL_REFDIV;
output	[2:0]	SP2HP_xPLL_VCO_Ctuning;
output	[2:0]	SP2HP_xPLL_buf_Itrim;
output		SP2HP_xPLL_lockdet_en;
output	[1:0]	SP2HP_xPLL_lockdet_period_sel;
output	[2:0]	SP2HP_xPLL_lockdet_ppm_sel1;
output	[2:0]	SP2HP_xPLL_lockdet_ppm_sel0;
output	[1:0]	SP2HP_xPLL_pdivSel;
output		SP2HP_xPLL_pwrdnB;
output		SP2HP_xPLL_resetB;
output		SP2HP_xPLL_selFourFive;
output		SP2HP_xRX3_busdivSel;
output		SP2HP_xRX3_pwrdnB;
output		SP2HP_xRX3_set_phase;
output		SP2HP_xRX3_slip_clk;
output		SP2HP_xRX3_syncRxToUsrclk;
output		SP2HP_xRX3_xrChicoOvrPh5to9;
output	[4:0]	SP2HP_xRX3_xrChicoOvrd;
output		SP2HP_xRX3_xrChicoOvrdEn;
output		SP2HP_xRX2_busdivSel;
output		SP2HP_xRX2_pwrdnB;
output		SP2HP_xRX2_set_phase;
output		SP2HP_xRX2_slip_clk;
output		SP2HP_xRX2_syncRxToUsrclk;
output		SP2HP_xRX2_xrChicoOvrPh5to9;
output	[4:0]	SP2HP_xRX2_xrChicoOvrd;
output		SP2HP_xRX2_xrChicoOvrdEn;
output		SP2HP_xRX1_busdivSel;
output		SP2HP_xRX1_pwrdnB;
output		SP2HP_xRX1_set_phase;
output		SP2HP_xRX1_slip_clk;
output		SP2HP_xRX1_syncRxToUsrclk;
output		SP2HP_xRX1_xrChicoOvrPh5to9;
output	[4:0]	SP2HP_xRX1_xrChicoOvrd;
output		SP2HP_xRX1_xrChicoOvrdEn;
output		SP2HP_xRX0_busdivSel;
output		SP2HP_xRX0_pwrdnB;
output		SP2HP_xRX0_set_phase;
output		SP2HP_xRX0_slip_clk;
output		SP2HP_xRX0_syncRxToUsrclk;
output		SP2HP_xRX0_xrChicoOvrPh5to9;
output	[4:0]	SP2HP_xRX0_xrChicoOvrd;
output		SP2HP_xRX0_xrChicoOvrdEn;
output	[1:0]	SP2HP_xRXAFE3_InCMTrim;
output		SP2HP_xRXAFE3_rcvShuntEn;
output		SP2HP_xRXAFE3_rcvVssTermEn;
output		SP2HP_xRXAFE3_rcvVttTermEn;
output		SP2HP_xRXAFE3_termRes50En;
output	[1:0]	SP2HP_xRXAFE2_InCMTrim;
output		SP2HP_xRXAFE2_rcvShuntEn;
output		SP2HP_xRXAFE2_rcvVssTermEn;
output		SP2HP_xRXAFE2_rcvVttTermEn;
output		SP2HP_xRXAFE2_termRes50En;
output	[1:0]	SP2HP_xRXAFE1_InCMTrim;
output		SP2HP_xRXAFE1_rcvShuntEn;
output		SP2HP_xRXAFE1_rcvVssTermEn;
output		SP2HP_xRXAFE1_rcvVttTermEn;
output		SP2HP_xRXAFE1_termRes50En;
output	[1:0]	SP2HP_xRXAFE0_InCMTrim;
output		SP2HP_xRXAFE0_rcvShuntEn;
output		SP2HP_xRXAFE0_rcvVssTermEn;
output		SP2HP_xRXAFE0_rcvVttTermEn;
output		SP2HP_xRXAFE0_termRes50En;
output	[2:0]	SP2HP_xRXSquelch3_noSigLevel;
output		SP2HP_xRXSquelch3_pwrdnB;
output	[2:0]	SP2HP_xRXSquelch2_noSigLevel;
output		SP2HP_xRXSquelch2_pwrdnB;
output	[2:0]	SP2HP_xRXSquelch1_noSigLevel;
output		SP2HP_xRXSquelch1_pwrdnB;
output	[2:0]	SP2HP_xRXSquelch0_noSigLevel;
output		SP2HP_xRXSquelch0_pwrdnB;
output	[2:0]	SP2HP_xResCal_Bg_offset;
output	[2:0]	SP2HP_xResCal_LPF_offset;
output		SP2HP_xResCal_MemCtrl;
output		SP2HP_xResCal_MemEn;
output	[4:0]	SP2HP_xResCal_MemRes_Bg;
output	[4:0]	SP2HP_xResCal_MemRes_LPF;
output	[4:0]	SP2HP_xResCal_MemRes_Rx;
output	[4:0]	SP2HP_xResCal_MemRes_Tx;
output		SP2HP_xResCal_ResBg_sel;
output		SP2HP_xResCal_ResLPF_sel;
output		SP2HP_xResCal_ResRx_sel;
output		SP2HP_xResCal_ResTx_sel;
output	[2:0]	SP2HP_xResCal_Rx_offset;
output	[2:0]	SP2HP_xResCal_Tx_offset;
output	[4:0]	SP2HP_xTOP_DivOOB;
output	[4:0]	SP2HP_xTOP_DivSSC;
output	[4:0]	SP2HP_xTOP_DivSYS;
output		SP2HP_xTOP_SYSClkSel;
output		SP2HP_xTX3_ACCCLK_ROTATEH;
output		SP2HP_xTX3_ACC_DIN_SEL;
output	[1:0]	SP2HP_xTX3_ACC_NSEL;
output	[7:0]	SP2HP_xTX3_ACC_OVERRIDE;
output		SP2HP_xTX3_ACC_OVERRIDE_EN;
output		SP2HP_xTX3_ACC_ROTATE;
output		SP2HP_xTX3_ACC_UPDNSW;
output		SP2HP_xTX3_Clk_pwrdnB;
output	[2:0]	SP2HP_xTX3_DrvPostCursor;
output	[2:0]	SP2HP_xTX3_DrvPreCursor;
output		SP2HP_xTX3_Drv_pwrdnB;
output	[2:0]	SP2HP_xTX3_Drvbiastrim;
output	[3:0]	SP2HP_xTX3_Drvswing;
output	[2:0]	SP2HP_xTX3_PI_captrim;
output		SP2HP_xTX3_PI_pwrdnB;
output	[1:0]	SP2HP_xTX3_PIbiasTrim;
output		SP2HP_xTX3_Resl_En;
output		SP2HP_xTX3_SSC_EN;
output	[8:0]	SP2HP_xTX3_SSC_OVERRIDE;
output		SP2HP_xTX3_SSC_OVERRIDE_EN;
output	[4:0]	SP2HP_xTX3_SSC_TSEL;
output		SP2HP_xTX3_Ser_pwrdnB;
output	[2:0]	SP2HP_xTX3_Serbiastrim;
output	[3:0]	SP2HP_xTX3_Vreftrim;
output		SP2HP_xTX3_activepkEn;
output		SP2HP_xTX3_busdivSel;
output		SP2HP_xTX3_chico_cksel;
output		SP2HP_xTX3_chico_pwrdnB;
output	[2:0]	SP2HP_xTX3_ctune;
output	[1:0]	SP2HP_xTX3_dccbiastrim;
output	[1:0]	SP2HP_xTX3_dccerrtrim;
output		SP2HP_xTX3_dccfix;
output	[2:0]	SP2HP_xTX3_gmtune;
output		SP2HP_xTX3_ovsdivEn;
output	[1:0]	SP2HP_xTX3_pdivSel;
output		SP2HP_xTX3_pwrdnB;
output		SP2HP_xTX3_selFourFive;
output		SP2HP_xTX3_sendidle;
output		SP2HP_xTX3_syncTxToUsrclk;
output		SP2HP_xTX3_tdccEn;
output		SP2HP_xTX3_tdccovrd;
output		SP2HP_xTX2_ACCCLK_ROTATEH;
output		SP2HP_xTX2_ACC_DIN_SEL;
output	[1:0]	SP2HP_xTX2_ACC_NSEL;
output	[7:0]	SP2HP_xTX2_ACC_OVERRIDE;
output		SP2HP_xTX2_ACC_OVERRIDE_EN;
output		SP2HP_xTX2_ACC_ROTATE;
output		SP2HP_xTX2_ACC_UPDNSW;
output		SP2HP_xTX2_Clk_pwrdnB;
output	[2:0]	SP2HP_xTX2_DrvPostCursor;
output	[2:0]	SP2HP_xTX2_DrvPreCursor;
output		SP2HP_xTX2_Drv_pwrdnB;
output	[2:0]	SP2HP_xTX2_Drvbiastrim;
output	[3:0]	SP2HP_xTX2_Drvswing;
output	[2:0]	SP2HP_xTX2_PI_captrim;
output		SP2HP_xTX2_PI_pwrdnB;
output	[1:0]	SP2HP_xTX2_PIbiasTrim;
output		SP2HP_xTX2_Resl_En;
output		SP2HP_xTX2_SSC_EN;
output	[8:0]	SP2HP_xTX2_SSC_OVERRIDE;
output		SP2HP_xTX2_SSC_OVERRIDE_EN;
output	[4:0]	SP2HP_xTX2_SSC_TSEL;
output		SP2HP_xTX2_Ser_pwrdnB;
output	[2:0]	SP2HP_xTX2_Serbiastrim;
output	[3:0]	SP2HP_xTX2_Vreftrim;
output		SP2HP_xTX2_activepkEn;
output		SP2HP_xTX2_busdivSel;
output		SP2HP_xTX2_chico_cksel;
output		SP2HP_xTX2_chico_pwrdnB;
output	[2:0]	SP2HP_xTX2_ctune;
output	[1:0]	SP2HP_xTX2_dccbiastrim;
output	[1:0]	SP2HP_xTX2_dccerrtrim;
output		SP2HP_xTX2_dccfix;
output	[2:0]	SP2HP_xTX2_gmtune;
output		SP2HP_xTX2_ovsdivEn;
output	[1:0]	SP2HP_xTX2_pdivSel;
output		SP2HP_xTX2_pwrdnB;
output		SP2HP_xTX2_selFourFive;
output		SP2HP_xTX2_sendidle;
output		SP2HP_xTX2_syncTxToUsrclk;
output		SP2HP_xTX2_tdccEn;
output		SP2HP_xTX2_tdccovrd;
output		SP2HP_xTX1_ACCCLK_ROTATEH;
output		SP2HP_xTX1_ACC_DIN_SEL;
output	[1:0]	SP2HP_xTX1_ACC_NSEL;
output	[7:0]	SP2HP_xTX1_ACC_OVERRIDE;
output		SP2HP_xTX1_ACC_OVERRIDE_EN;
output		SP2HP_xTX1_ACC_ROTATE;
output		SP2HP_xTX1_ACC_UPDNSW;
output		SP2HP_xTX1_Clk_pwrdnB;
output	[2:0]	SP2HP_xTX1_DrvPostCursor;
output	[2:0]	SP2HP_xTX1_DrvPreCursor;
output		SP2HP_xTX1_Drv_pwrdnB;
output	[2:0]	SP2HP_xTX1_Drvbiastrim;
output	[3:0]	SP2HP_xTX1_Drvswing;
output	[2:0]	SP2HP_xTX1_PI_captrim;
output		SP2HP_xTX1_PI_pwrdnB;
output	[1:0]	SP2HP_xTX1_PIbiasTrim;
output		SP2HP_xTX1_Resl_En;
output		SP2HP_xTX1_SSC_EN;
output	[8:0]	SP2HP_xTX1_SSC_OVERRIDE;
output		SP2HP_xTX1_SSC_OVERRIDE_EN;
output	[4:0]	SP2HP_xTX1_SSC_TSEL;
output		SP2HP_xTX1_Ser_pwrdnB;
output	[2:0]	SP2HP_xTX1_Serbiastrim;
output	[3:0]	SP2HP_xTX1_Vreftrim;
output		SP2HP_xTX1_activepkEn;
output		SP2HP_xTX1_busdivSel;
output		SP2HP_xTX1_chico_cksel;
output		SP2HP_xTX1_chico_pwrdnB;
output	[2:0]	SP2HP_xTX1_ctune;
output	[1:0]	SP2HP_xTX1_dccbiastrim;
output	[1:0]	SP2HP_xTX1_dccerrtrim;
output		SP2HP_xTX1_dccfix;
output	[2:0]	SP2HP_xTX1_gmtune;
output		SP2HP_xTX1_ovsdivEn;
output	[1:0]	SP2HP_xTX1_pdivSel;
output		SP2HP_xTX1_pwrdnB;
output		SP2HP_xTX1_selFourFive;
output		SP2HP_xTX1_sendidle;
output		SP2HP_xTX1_syncTxToUsrclk;
output		SP2HP_xTX1_tdccEn;
output		SP2HP_xTX1_tdccovrd;
output		SP2HP_xTX0_ACCCLK_ROTATEH;
output		SP2HP_xTX0_ACC_DIN_SEL;
output	[1:0]	SP2HP_xTX0_ACC_NSEL;
output	[7:0]	SP2HP_xTX0_ACC_OVERRIDE;
output		SP2HP_xTX0_ACC_OVERRIDE_EN;
output		SP2HP_xTX0_ACC_ROTATE;
output		SP2HP_xTX0_ACC_UPDNSW;
output		SP2HP_xTX0_Clk_pwrdnB;
output	[2:0]	SP2HP_xTX0_DrvPostCursor;
output	[2:0]	SP2HP_xTX0_DrvPreCursor;
output		SP2HP_xTX0_Drv_pwrdnB;
output	[2:0]	SP2HP_xTX0_Drvbiastrim;
output	[3:0]	SP2HP_xTX0_Drvswing;
output	[2:0]	SP2HP_xTX0_PI_captrim;
output		SP2HP_xTX0_PI_pwrdnB;
output	[1:0]	SP2HP_xTX0_PIbiasTrim;
output		SP2HP_xTX0_Resl_En;
output		SP2HP_xTX0_SSC_EN;
output	[8:0]	SP2HP_xTX0_SSC_OVERRIDE;
output		SP2HP_xTX0_SSC_OVERRIDE_EN;
output	[4:0]	SP2HP_xTX0_SSC_TSEL;
output		SP2HP_xTX0_Ser_pwrdnB;
output	[2:0]	SP2HP_xTX0_Serbiastrim;
output	[3:0]	SP2HP_xTX0_Vreftrim;
output		SP2HP_xTX0_activepkEn;
output		SP2HP_xTX0_busdivSel;
output		SP2HP_xTX0_chico_cksel;
output		SP2HP_xTX0_chico_pwrdnB;
output	[2:0]	SP2HP_xTX0_ctune;
output	[1:0]	SP2HP_xTX0_dccbiastrim;
output	[1:0]	SP2HP_xTX0_dccerrtrim;
output		SP2HP_xTX0_dccfix;
output	[2:0]	SP2HP_xTX0_gmtune;
output		SP2HP_xTX0_ovsdivEn;
output	[1:0]	SP2HP_xTX0_pdivSel;
output		SP2HP_xTX0_pwrdnB;
output		SP2HP_xTX0_selFourFive;
output		SP2HP_xTX0_sendidle;
output		SP2HP_xTX0_syncTxToUsrclk;
output		SP2HP_xTX0_tdccEn;
output		SP2HP_xTX0_tdccovrd;
output		SP2HP_xTX_SSC_Align;
output		SP2LP_pipe0_phystatus;
output	[2:0]	app_parity_errs;
output	[0:0]	aux_pm_en;
output		cfg_2nd_reset;
output	[7:0]	cfg_2ndbus_num;
output	[4:0]	cfg_aer_int_msg_num;
output	[0:0]	cfg_aer_rc_err_int;
output	[0:0]	cfg_aer_rc_err_msi;
output	[1:0]	cfg_atten_ind;
output	[31:0]	cfg_bar5_limit;
output	[31:0]	cfg_bar5_start;
output	[63:0]	cfg_bar4_limit;
output	[63:0]	cfg_bar4_start;
output	[31:0]	cfg_bar3_limit;
output	[31:0]	cfg_bar3_start;
output	[63:0]	cfg_bar2_limit;
output	[63:0]	cfg_bar2_start;
output	[31:0]	cfg_bar1_limit;
output	[31:0]	cfg_bar1_start;
output	[63:0]	cfg_bar0_limit;
output	[63:0]	cfg_bar0_start;
output	[0:0]	cfg_bus_master_en;
output		cfg_bw_mgt_int;
output	[0:0]	cfg_eml_control;
output	[31:0]	cfg_exp_rom_limit;
output	[31:0]	cfg_exp_rom_start;
output	[0:0]	cfg_int_disable;
output		cfg_link_auto_bw_int;
output	[2:0]	cfg_max_payload_size;
output	[2:0]	cfg_max_rd_req_size;
output	[0:0]	cfg_mem_space_en;
output	[0:0]	cfg_msi_64;
output	[63:0]	cfg_msi_addr;
output	[15:0]	cfg_msi_data;
output	[0:0]	cfg_msi_en;
output	[31:0]	cfg_msi_mask;
output	[2:0]	cfg_multi_msi_en;
output	[0:0]	cfg_no_snoop_en;
output	[4:0]	cfg_pbus_dev_num;
output	[7:0]	cfg_pbus_num;
output	[4:0]	cfg_pcie_cap_int_msg_num;
output	[0:0]	cfg_pm_no_soft_rst;
output	[0:0]	cfg_pme_int;
output	[0:0]	cfg_pme_msi;
output	[0:0]	cfg_pwr_ctrler_ctrl;
output	[1:0]	cfg_pwr_ind;
output	[0:0]	cfg_rcb;
output	[0:0]	cfg_relax_order_en;
output	[0:0]	cfg_send_cor_err;
output	[0:0]	cfg_send_f_err;
output	[0:0]	cfg_send_nf_err;
output	[7:0]	cfg_subbus_num;
output	[0:0]	cfg_sys_err_rc;
output		clk_req_n;
output	[63:0]	cxpl_debug_info;
output	[15:0]	cxpl_debug_info_ei;
output	[801:0]	diag_status_bus;
output		en_aux_clk_g;
output	[0:0]	hp_int;
output	[0:0]	hp_msi;
output	[0:0]	hp_pme;
output		lbc_dbi_ack;
output	[31:0]	lbc_dbi_dout;
output	[15:0]	lbc_ext_addr;
output	[2:0]	lbc_ext_bar_num;
output	[0:0]	lbc_ext_cs;
output	[31:0]	lbc_ext_dout;
output		lbc_ext_io_access;
output		lbc_ext_rom_access;
output	[3:0]	lbc_ext_wr;
output		link_req_rst_not;
output		mac_phy_rate;
output	[3:0]	mac_phy_rxstandby;
output	[2:0]	pm_curnt_state;
output	[2:0]	pm_dstate;
output		pm_linkst_in_l2;
output		pm_linkst_in_l1;
output		pm_linkst_in_l0s;
output		pm_linkst_l2_exit;
output	[0:0]	pm_pme_en;
output		pm_req_core_rst;
output		pm_req_non_sticky_rst;
output		pm_req_phy_rst;
output		pm_req_sticky_rst;
output		pm_sel_aux_clk;
output	[0:0]	pm_status;
output		pm_xtlh_block_tlp;
output	[63:0]	radm_bypass_addr;
output	[1:0]	radm_bypass_attr;
output	[0:0]	radm_bypass_bcm;
output	[11:0]	radm_bypass_byte_cnt;
output	[15:0]	radm_bypass_cmpltr_id;
output	[0:0]	radm_bypass_cpl_last;
output	[2:0]	radm_bypass_cpl_status;
output	[127:0]	radm_bypass_data;
output	[0:0]	radm_bypass_dllp_abort;
output	[0:0]	radm_bypass_dv;
output	[9:0]	radm_bypass_dw_len;
output	[3:0]	radm_bypass_dwen;
output	[0:0]	radm_bypass_ecrc_err;
output	[0:0]	radm_bypass_eot;
output	[3:0]	radm_bypass_first_be;
output	[1:0]	radm_bypass_fmt;
output	[2:0]	radm_bypass_func_num;
output	[0:0]	radm_bypass_hv;
output	[2:0]	radm_bypass_in_membar_range;
output	[0:0]	radm_bypass_io_req_in_range;
output	[3:0]	radm_bypass_last_be;
output	[0:0]	radm_bypass_poisoned;
output	[15:0]	radm_bypass_reqid;
output	[0:0]	radm_bypass_rom_in_range;
output	[7:0]	radm_bypass_tag;
output	[2:0]	radm_bypass_tc;
output	[0:0]	radm_bypass_td;
output	[0:0]	radm_bypass_tlp_abort;
output	[4:0]	radm_bypass_type;
output		radm_correctable_err;
output		radm_cpl_timeout;
output		radm_fatal_err;
output	[11:0]	radm_grant_tlp_type;
output		radm_inta_asserted;
output		radm_inta_deasserted;
output		radm_intb_asserted;
output		radm_intb_deasserted;
output		radm_intc_asserted;
output		radm_intc_deasserted;
output		radm_intd_asserted;
output		radm_intd_deasserted;
output	[63:0]	radm_msg_payload;
output	[15:0]	radm_msg_req_id;
output		radm_msg_unlock;
output		radm_nonfatal_err;
output	[0:0]	radm_pm_pme;
output		radm_pm_to_ack;
output		radm_pm_turnoff;
output	[3:0]	radm_q_not_empty;
output	[3:0]	radm_qoverflow;
output	[1:0]	radm_timeout_cpl_attr;
output	[11:0]	radm_timeout_cpl_len;
output	[7:0]	radm_timeout_cpl_tag;
output	[2:0]	radm_timeout_cpl_tc;
output	[2:0]	radm_timeout_func_num;
output	[63:0]	radm_trgt1_addr;
output	[1:0]	radm_trgt1_attr;
output		radm_trgt1_bcm;
output	[11:0]	radm_trgt1_byte_cnt;
output	[15:0]	radm_trgt1_cmpltr_id;
output		radm_trgt1_cpl_last;
output	[2:0]	radm_trgt1_cpl_status;
output	[127:0]	radm_trgt1_data;
output		radm_trgt1_dllp_abort;
output		radm_trgt1_dv;
output	[9:0]	radm_trgt1_dw_len;
output	[3:0]	radm_trgt1_dwen;
output		radm_trgt1_ecrc_err;
output		radm_trgt1_eot;
output	[3:0]	radm_trgt1_first_be;
output	[1:0]	radm_trgt1_fmt;
output	[2:0]	radm_trgt1_func_num;
output		radm_trgt1_hv;
output	[2:0]	radm_trgt1_in_membar_range;
output		radm_trgt1_io_req_in_range;
output	[3:0]	radm_trgt1_last_be;
output		radm_trgt1_mem_type;
output		radm_trgt1_poisoned;
output	[15:0]	radm_trgt1_reqid;
output		radm_trgt1_rom_in_range;
output	[7:0]	radm_trgt1_tag;
output	[2:0]	radm_trgt1_tc;
output		radm_trgt1_td;
output		radm_trgt1_tlp_abort;
output	[4:0]	radm_trgt1_type;
output	[0:0]	radm_vendor_msg;
output		rdlh_link_up;
output		routing_pipe_glue_rstn;
output	[63:0]	rtlh_rfc_data;
output	[1:0]	rtlh_rfc_upd;
output		smlh_link_up;
output	[5:0]	smlh_ltssm_state;
output		smlh_req_rst_not;
output		training_rst_n;
output		trgt_cpl_timeout;
output		trgt_lookup_empty;
output	[7:0]	trgt_lookup_id;
output	[1:0]	trgt_timeout_cpl_attr;
output	[2:0]	trgt_timeout_cpl_func_num;
output	[11:0]	trgt_timeout_cpl_len;
output	[2:0]	trgt_timeout_cpl_tc;
output	[7:0]	trgt_timeout_lookup_id;
output		ven_msg_grant;
output		ven_msi_grant;
output		wake;
output		xadm_client1_halt;
output		xadm_client0_halt;
output	[47:0]	xadm_cpld_cdts;
output	[31:0]	xadm_cplh_cdts;
output	[47:0]	xadm_npd_cdts;
output	[31:0]	xadm_nph_cdts;
output	[47:0]	xadm_pd_cdts;
output	[31:0]	xadm_ph_cdts;
input		HP2SP_L3RxCALDetected;
input		HP2SP_L3RxGearboxIsSync;
input		HP2SP_L3RxOOBCOMINITDet;
input		HP2SP_L3RxOOBCOMSASDet;
input		HP2SP_L3RxOOBCOMWAKEDet;
input		HP2SP_L3RxOOBElecIdle;
input		HP2SP_L3RxOvrsmplErr;
input		HP2SP_L3RxPIPEPHYStatusRxDet;
input		HP2SP_L3RxPIPERxDetected;
input	[15:0]	HP2SP_L3RxPRBSErrCnt;
input	[15:0]	HP2SP_L3RxPRBSZeroCnt;
input		HP2SP_L3RxRecClk;
input		HP2SP_L3RxRecClk2;
input	[1:0]	HP2SP_L3RxSyncState;
input	[7:0]	HP2SP_L3RxUsr8B10BDispErr;
input	[11:0]	HP2SP_L3RxUsr8B10BEBCorCnt;
input	[11:0]	HP2SP_L3RxUsr8B10BEBStat;
input	[7:0]	HP2SP_L3RxUsr8B10BIsComma;
input	[7:0]	HP2SP_L3RxUsr8B10BIsK;
input	[7:0]	HP2SP_L3RxUsr8B10BNotInTable;
input	[7:0]	HP2SP_L3RxUsr8B10BRunDisp;
input		HP2SP_L3RxUsr8B10BValid;
input	[79:0]	HP2SP_L3RxUsrData;
input		HP2SP_L3RxUsrDataValid;
input	[2:0]	HP2SP_L3RxUsrGBHeader;
input		HP2SP_L3RxUsrGBHeaderValid;
input		HP2SP_L3RxUsrGBStartSeq;
input	[2:0]	HP2SP_L3TxBufStatus;
input		HP2SP_L3TxOutClk;
input		HP2SP_L3TxOutClk2;
input		HP2SP_L3TxSATAOOBComFinish;
input		HP2SP_L3TxUsrGBReady;
input		HP2SP_L2RxCALDetected;
input		HP2SP_L2RxGearboxIsSync;
input		HP2SP_L2RxOOBCOMINITDet;
input		HP2SP_L2RxOOBCOMSASDet;
input		HP2SP_L2RxOOBCOMWAKEDet;
input		HP2SP_L2RxOOBElecIdle;
input		HP2SP_L2RxOvrsmplErr;
input		HP2SP_L2RxPIPEPHYStatusRxDet;
input		HP2SP_L2RxPIPERxDetected;
input	[15:0]	HP2SP_L2RxPRBSErrCnt;
input	[15:0]	HP2SP_L2RxPRBSZeroCnt;
input		HP2SP_L2RxRecClk;
input		HP2SP_L2RxRecClk2;
input	[1:0]	HP2SP_L2RxSyncState;
input	[7:0]	HP2SP_L2RxUsr8B10BDispErr;
input	[11:0]	HP2SP_L2RxUsr8B10BEBCorCnt;
input	[11:0]	HP2SP_L2RxUsr8B10BEBStat;
input	[7:0]	HP2SP_L2RxUsr8B10BIsComma;
input	[7:0]	HP2SP_L2RxUsr8B10BIsK;
input	[7:0]	HP2SP_L2RxUsr8B10BNotInTable;
input	[7:0]	HP2SP_L2RxUsr8B10BRunDisp;
input		HP2SP_L2RxUsr8B10BValid;
input	[79:0]	HP2SP_L2RxUsrData;
input		HP2SP_L2RxUsrDataValid;
input	[2:0]	HP2SP_L2RxUsrGBHeader;
input		HP2SP_L2RxUsrGBHeaderValid;
input		HP2SP_L2RxUsrGBStartSeq;
input	[2:0]	HP2SP_L2TxBufStatus;
input		HP2SP_L2TxOutClk;
input		HP2SP_L2TxOutClk2;
input		HP2SP_L2TxSATAOOBComFinish;
input		HP2SP_L2TxUsrGBReady;
input		HP2SP_L1RxCALDetected;
input		HP2SP_L1RxGearboxIsSync;
input		HP2SP_L1RxOOBCOMINITDet;
input		HP2SP_L1RxOOBCOMSASDet;
input		HP2SP_L1RxOOBCOMWAKEDet;
input		HP2SP_L1RxOOBElecIdle;
input		HP2SP_L1RxOvrsmplErr;
input		HP2SP_L1RxPIPEPHYStatusRxDet;
input		HP2SP_L1RxPIPERxDetected;
input	[15:0]	HP2SP_L1RxPRBSErrCnt;
input	[15:0]	HP2SP_L1RxPRBSZeroCnt;
input		HP2SP_L1RxRecClk;
input		HP2SP_L1RxRecClk2;
input	[1:0]	HP2SP_L1RxSyncState;
input	[7:0]	HP2SP_L1RxUsr8B10BDispErr;
input	[11:0]	HP2SP_L1RxUsr8B10BEBCorCnt;
input	[11:0]	HP2SP_L1RxUsr8B10BEBStat;
input	[7:0]	HP2SP_L1RxUsr8B10BIsComma;
input	[7:0]	HP2SP_L1RxUsr8B10BIsK;
input	[7:0]	HP2SP_L1RxUsr8B10BNotInTable;
input	[7:0]	HP2SP_L1RxUsr8B10BRunDisp;
input		HP2SP_L1RxUsr8B10BValid;
input	[79:0]	HP2SP_L1RxUsrData;
input		HP2SP_L1RxUsrDataValid;
input	[2:0]	HP2SP_L1RxUsrGBHeader;
input		HP2SP_L1RxUsrGBHeaderValid;
input		HP2SP_L1RxUsrGBStartSeq;
input	[2:0]	HP2SP_L1TxBufStatus;
input		HP2SP_L1TxOutClk;
input		HP2SP_L1TxOutClk2;
input		HP2SP_L1TxSATAOOBComFinish;
input		HP2SP_L1TxUsrGBReady;
input		HP2SP_L0RxCALDetected;
input		HP2SP_L0RxGearboxIsSync;
input		HP2SP_L0RxOOBCOMINITDet;
input		HP2SP_L0RxOOBCOMSASDet;
input		HP2SP_L0RxOOBCOMWAKEDet;
input		HP2SP_L0RxOOBElecIdle;
input		HP2SP_L0RxOvrsmplErr;
input		HP2SP_L0RxPIPEPHYStatusRxDet;
input		HP2SP_L0RxPIPERxDetected;
input	[15:0]	HP2SP_L0RxPRBSErrCnt;
input	[15:0]	HP2SP_L0RxPRBSZeroCnt;
input		HP2SP_L0RxRecClk;
input		HP2SP_L0RxRecClk2;
input	[1:0]	HP2SP_L0RxSyncState;
input	[7:0]	HP2SP_L0RxUsr8B10BDispErr;
input	[11:0]	HP2SP_L0RxUsr8B10BEBCorCnt;
input	[11:0]	HP2SP_L0RxUsr8B10BEBStat;
input	[7:0]	HP2SP_L0RxUsr8B10BIsComma;
input	[7:0]	HP2SP_L0RxUsr8B10BIsK;
input	[7:0]	HP2SP_L0RxUsr8B10BNotInTable;
input	[7:0]	HP2SP_L0RxUsr8B10BRunDisp;
input		HP2SP_L0RxUsr8B10BValid;
input	[79:0]	HP2SP_L0RxUsrData;
input		HP2SP_L0RxUsrDataValid;
input	[2:0]	HP2SP_L0RxUsrGBHeader;
input		HP2SP_L0RxUsrGBHeaderValid;
input		HP2SP_L0RxUsrGBStartSeq;
input	[2:0]	HP2SP_L0TxBufStatus;
input		HP2SP_L0TxOutClk;
input		HP2SP_L0TxOutClk2;
input		HP2SP_L0TxSATAOOBComFinish;
input		HP2SP_L0TxUsrGBReady;
input		HP2SP_PIPEPhyStatusForce;
input		HP2SP_PIPEPhyStatusSoft;
input		HP2SP_PowerOnDone;
input		HP2SP_RxLDuAlignAcqr;
input		HP2SP_SysClk;
input		HP2SP_xPLL_DivClk;
input		app_clk_req_n;
input	[3:0]	app_cpld_ca;
input	[3:0]	app_cplh_ca;
input		app_err_advisory;
input	[11:0]	app_err_bus;
input	[2:0]	app_err_func_num;
input	[127:0]	app_hdr_log;
input		app_hdr_valid;
input		app_init_rst;
input		app_ltssm_enable;
input	[3:0]	app_npd_ca;
input	[3:0]	app_nph_ca;
input	[3:0]	app_pd_ca;
input	[3:0]	app_ph_ca;
input		app_ready_entr_l23;
input		app_req_entr_l1;
input		app_req_exit_l1;
input		app_req_retry_en;
input		app_unlock_msg;
input		app_xfer_pending;
input	[0:0]	apps_pm_xmt_pme;
input		apps_pm_xmt_turnoff;
input		aux_clk;
input		aux_clk_active;
input		aux_clk_g;
input	[31:0]	cfg_msi_pending;
input		client1_addr_align_en;
input		client1_cpl_bcm;
input	[11:0]	client1_cpl_byte_cnt;
input	[7:0]	client1_cpl_lookup_id;
input	[2:0]	client1_cpl_status;
input	[15:0]	client1_remote_req_id;
input	[65:0]	client1_tlp_addr;
input	[1:0]	client1_tlp_attr;
input		client1_tlp_bad_eot;
input	[7:0]	client1_tlp_byte_en;
input	[12:0]	client1_tlp_byte_len;
input	[131:0]	client1_tlp_data;
input		client1_tlp_dv;
input		client1_tlp_eot;
input		client1_tlp_ep;
input	[1:0]	client1_tlp_fmt;
input	[2:0]	client1_tlp_func_num;
input		client1_tlp_hv;
input	[2:0]	client1_tlp_tc;
input		client1_tlp_td;
input	[7:0]	client1_tlp_tid;
input	[4:0]	client1_tlp_type;
input		client0_addr_align_en;
input		client0_cpl_bcm;
input	[11:0]	client0_cpl_byte_cnt;
input	[7:0]	client0_cpl_lookup_id;
input	[2:0]	client0_cpl_status;
input	[15:0]	client0_remote_req_id;
input	[65:0]	client0_tlp_addr;
input	[1:0]	client0_tlp_attr;
input		client0_tlp_bad_eot;
input	[7:0]	client0_tlp_byte_en;
input	[12:0]	client0_tlp_byte_len;
input	[131:0]	client0_tlp_data;
input		client0_tlp_dv;
input		client0_tlp_eot;
input		client0_tlp_ep;
input	[1:0]	client0_tlp_fmt;
input	[2:0]	client0_tlp_func_num;
input		client0_tlp_hv;
input	[2:0]	client0_tlp_tc;
input		client0_tlp_td;
input	[7:0]	client0_tlp_tid;
input	[4:0]	client0_tlp_type;
input		core_clk;
input		core_clk_ug;
input		core_rst_n;
input		dbg_pba;
input		dbg_table;
input	[31:0]	fp_dbi_addr;
input	[2:0]	fp_dbi_bar_num;
input		fp_dbi_cs;
input		fp_dbi_cs2;
input	[31:0]	fp_dbi_din;
input	[2:0]	fp_dbi_func_num;
input		fp_dbi_io_access;
input		fp_dbi_rom_access;
input	[3:0]	fp_dbi_wr;
input	[31:0]	ccb_dbi_addr;
input	[2:0]	ccb_dbi_bar_num;
input		ccb_dbi_cs;
input		ccb_dbi_cs2;
input	[31:0]	ccb_dbi_din;
input	[2:0]	ccb_dbi_func_num;
input		ccb_dbi_io_access;
input		ccb_dbi_rom_access;
input	[3:0]	ccb_dbi_wr;
input		ccb_lbc_dbi_ack;
input	[31:0]	ccb_lbc_dbi_dout;
output		cbi_pbus_gnt;
output	[31:0]	cbi_pbus_rdata;
input		clk_p;
input		rst_p_n;
input	[15:0]	cbi_pbus_addr;
input		cbi_pbus_write;
input		cbi_pbus_req;
input	[31:0]	cbi_pbus_wdata;
input	[3:0]	device_type;
input	[2:0]	diag_ctrl_bus;
input	[0:0]	ext_lbc_ack;
input	[31:0]	ext_lbc_din;
input		fp2HP_pcs_usr_resetB;
input		fp2LP_pipe_glue_rstn;
input		non_sticky_rst_n;
input	[0:0]	outband_pwrup_cmd;
input		perst_n;
input		phy_clk_req_n;
input		pipe_clk;
input		pipe_glue_rstn;
input		pipe_rst_n;
input		pwr_rst_n;
input		rx_lane_flip_en;
input		squelch_rst_n;
input		sticky_rst_n;
input	[0:0]	sys_atten_button_pressed;
input		sys_aux_pwr_det;
input	[0:0]	sys_cmd_cpled_int;
input	[0:0]	sys_eml_interlock_engaged;
input	[0:0]	sys_int;
input	[0:0]	sys_mrl_sensor_chged;
input	[0:0]	sys_mrl_sensor_state;
input	[0:0]	sys_pre_det_chged;
input	[0:0]	sys_pre_det_state;
input	[0:0]	sys_pwr_fault_det;
input		trgt1_radm_halt;
input	[11:0]	trgt1_radm_pkt_halt;
input		tx_lane_flip_en;
input	[1:0]	ven_msg_attr;
input	[7:0]	ven_msg_code;
input	[63:0]	ven_msg_data;
input		ven_msg_ep;
input	[1:0]	ven_msg_fmt;
input	[2:0]	ven_msg_func_num;
input	[9:0]	ven_msg_len;
input		ven_msg_req;
input	[7:0]	ven_msg_tag;
input	[2:0]	ven_msg_tc;
input		ven_msg_td;
input	[4:0]	ven_msg_type;
input	[2:0]	ven_msi_func_num;
input		ven_msi_req;
input	[2:0]	ven_msi_tc;
input	[4:0]	ven_msi_vector;

parameter cfg_dbimux_ccb_fp  = 1'b0;  //0: ccb, 1: FP
parameter pcie_iso_en = 1'b0;
parameter cfg_reg_cbi = 8'b0;

endmodule

// VPERL: GENERATED_BEG

module phy_wrapper (
	ahb_hrdata_o,
	ahb_hready_o,
	ahb_hresp_o,
	dram_dfi_ctrlupd_ack,
	dram_dfi_ecc_rddata_w1,
	dram_dfi_ecc_rddata_w0,
	dram_dfi_init_complete,
	dram_dfi_rddata_valid_w1,
	dram_dfi_rddata_valid_w0,
	dram_dfi_rddata_w1,
	dram_dfi_rddata_w0,
	dram_dfi_rdlvl_gate_mode,
	dram_dfi_rdlvl_mode,
	dram_dfi_rdlvl_resp,
	dram_dfi_wrlvl_mode,
	dram_dfi_wrlvl_resp,
	fp_dfi_ctrlupd_ack,
	fp_dfi_ecc_rddata_valid_w1,
	fp_dfi_ecc_rddata_valid_w0,
	fp_dfi_ecc_rddata_w1,
	fp_dfi_ecc_rddata_w0,
	fp_dfi_init_complete,
	fp_dfi_rddata_valid_w1,
	fp_dfi_rddata_valid_w0,
	fp_dfi_rddata_w1,
	fp_dfi_rddata_w0,
	fp_dfi_rdlvl_gate_mode,
	fp_dfi_rdlvl_mode,
	fp_dfi_rdlvl_resp,
	fp_dfi_wrlvl_mode,
	fp_dfi_wrlvl_resp,
	iodc_jtag_ddr_addr_c,
	iodc_jtag_ddr_bank_c,
	iodc_jtag_ddr_cas_n_c,
	iodc_jtag_ddr_cke_c,
	iodc_jtag_ddr_clk_c,
	iodc_jtag_ddr_cs_n_c,
	iodc_jtag_ddr_dm_c,
	iodc_jtag_ddr_dq_c,
	iodc_jtag_ddr_dqs_c,
	iodc_jtag_ddr_ecc_dm_c,
	iodc_jtag_ddr_ecc_dq_c,
	iodc_jtag_ddr_ecc_dqs_c,
	iodc_jtag_ddr_odt_c,
	iodc_jtag_ddr_par_c,
	iodc_jtag_ddr_ras_n_c,
	iodc_jtag_ddr_reset_n_c,
	iodc_jtag_ddr_we_n_c,
//	phy_scan_out_d2f,
//	phy_scan_out_d2r,
//	phy_scan_out_x2f,
//	phy_scan_out_x2r,
	ro_ddr23phy_reg,
	ahb_haddr_i,
	ahb_hburst_i,
	ahb_hclk,
	ahb_hready_i,
	ahb_hresetn,
	ahb_hsel_i,
	ahb_hsize_i,
	ahb_htrans_i,
	ahb_hwdata_i,
	ahb_hwrite_i,
	bypasspll_mc_clk_x4,
//	dfi_sphy_sel,
	dram_dfi_addr_p1,
	dram_dfi_addr_p0,
	dram_dfi_bank_p1,
	dram_dfi_bank_p0,
	dram_dfi_cas_n_p1,
	dram_dfi_cas_n_p0,
	dram_dfi_cke_p1,
	dram_dfi_cke_p0,
	dram_dfi_cs_n_duplicate_p1,
	dram_dfi_cs_n_duplicate_p0,
	dram_dfi_cs_n_p1,
	dram_dfi_cs_n_p0,
	dram_dfi_ctrlupd_req,
	dram_dfi_dram_clk_disable,
	dram_dfi_ecc_rddata_en_p1,
	dram_dfi_ecc_rddata_en_p0,
	dram_dfi_ecc_wrdata_en_p1,
	dram_dfi_ecc_wrdata_en_p0,
	dram_dfi_ecc_wrdata_p1,
	dram_dfi_ecc_wrdata_p0,
	dram_dfi_ecc_wrmask_p1,
	dram_dfi_ecc_wrmask_p0,
	dram_dfi_init_start,
	dram_dfi_ras_n_p1,
	dram_dfi_ras_n_p0,
	dram_dfi_rddata_en_p1,
	dram_dfi_rddata_en_p0,
	dram_dfi_rdlvl_delay,
	dram_dfi_rdlvl_delayn,
	dram_dfi_rdlvl_edge,
	dram_dfi_rdlvl_en,
	dram_dfi_rdlvl_gate_delay,
	dram_dfi_rdlvl_gate_en,
	dram_dfi_rdlvl_load,
	dram_dfi_reset_n_p1,
	dram_dfi_reset_n_p0,
	dram_dfi_we_n_p1,
	dram_dfi_we_n_p0,
	dram_dfi_wodt_p1,
	dram_dfi_wodt_p0,
	dram_dfi_wrdata_en_p1,
	dram_dfi_wrdata_en_p0,
	dram_dfi_wrdata_p1,
	dram_dfi_wrdata_p0,
	dram_dfi_wrlvl_delay,
	dram_dfi_wrlvl_en,
	dram_dfi_wrlvl_load,
	dram_dfi_wrlvl_strobe,
	dram_dfi_wrmask_p1,
	dram_dfi_wrmask_p0,
	fp_dfi_addr_p1,
	fp_dfi_addr_p0,
	fp_dfi_bank_p1,
	fp_dfi_bank_p0,
	fp_dfi_cas_n_p1,
	fp_dfi_cas_n_p0,
	fp_dfi_cke_p1,
	fp_dfi_cke_p0,
	fp_dfi_cs_n_duplicate_p1,
	fp_dfi_cs_n_duplicate_p0,
	fp_dfi_cs_n_p1,
	fp_dfi_cs_n_p0,
	fp_dfi_ctrlupd_req,
	fp_dfi_dram_clk_disable,
	fp_dfi_ecc_rddata_en_p1,
	fp_dfi_ecc_rddata_en_p0,
	fp_dfi_ecc_wrdata_en_p1,
	fp_dfi_ecc_wrdata_en_p0,
	fp_dfi_ecc_wrdata_p1,
	fp_dfi_ecc_wrdata_p0,
	fp_dfi_ecc_wrmask_p1,
	fp_dfi_ecc_wrmask_p0,
	fp_dfi_init_start,
	fp_dfi_ras_n_p1,
	fp_dfi_ras_n_p0,
	fp_dfi_rddata_en_p1,
	fp_dfi_rddata_en_p0,
	fp_dfi_rdlvl_delay,
	fp_dfi_rdlvl_delayn,
	fp_dfi_rdlvl_edge,
	fp_dfi_rdlvl_en,
	fp_dfi_rdlvl_gate_delay,
	fp_dfi_rdlvl_gate_en,
	fp_dfi_rdlvl_load,
	fp_dfi_reset_n_p1,
	fp_dfi_reset_n_p0,
	fp_dfi_we_n_p1,
	fp_dfi_we_n_p0,
	fp_dfi_wodt_p1,
	fp_dfi_wodt_p0,
	fp_dfi_wrdata_en_p1,
	fp_dfi_wrdata_en_p0,
	fp_dfi_wrdata_p1,
	fp_dfi_wrdata_p0,
	fp_dfi_wrlvl_delay,
	fp_dfi_wrlvl_en,
	fp_dfi_wrlvl_load,
	fp_dfi_wrlvl_strobe,
	fp_dfi_wrmask_p1,
	fp_dfi_wrmask_p0,
	iodc_jtag_ddr_addr_i,
	iodc_jtag_ddr_addr_oe_n,
//	iodc_jtag_ddr_addr_pd,
//	iodc_jtag_ddr_addr_pu,
	iodc_jtag_ddr_bank_i,
	iodc_jtag_ddr_bank_oe_n,
//	iodc_jtag_ddr_bank_pd,
//	iodc_jtag_ddr_bank_pu,
	iodc_jtag_ddr_cas_n_i,
	iodc_jtag_ddr_cas_n_oe_n,
//	iodc_jtag_ddr_cas_n_pd,
//	iodc_jtag_ddr_cas_n_pu,
	iodc_jtag_ddr_cke_i,
	iodc_jtag_ddr_cke_oe_n,
//	iodc_jtag_ddr_cke_pd,
//	iodc_jtag_ddr_cke_pu,
	iodc_jtag_ddr_clk_i,
	iodc_jtag_ddr_clk_oe_n,
//	iodc_jtag_ddr_clk_pd,
//	iodc_jtag_ddr_clk_pu,
	iodc_jtag_ddr_cs_n_i,
	iodc_jtag_ddr_cs_n_oe_n,
//	iodc_jtag_ddr_cs_n_pd,
//	iodc_jtag_ddr_cs_n_pu,
	iodc_jtag_ddr_dm_i,
	iodc_jtag_ddr_dm_oe_n,
//	iodc_jtag_ddr_dm_pd,
//	iodc_jtag_ddr_dm_pu,
	iodc_jtag_ddr_dq_i,
	iodc_jtag_ddr_dq_oe_n,
//	iodc_jtag_ddr_dq_pd,
//	iodc_jtag_ddr_dq_pu,
	iodc_jtag_ddr_dqs_i,
	iodc_jtag_ddr_dqs_oe_n,
//	iodc_jtag_ddr_dqs_pd,
//	iodc_jtag_ddr_dqs_pu,
	iodc_jtag_ddr_ecc_dm_i,
	iodc_jtag_ddr_ecc_dm_oe_n,
//	iodc_jtag_ddr_ecc_dm_pd,
//	iodc_jtag_ddr_ecc_dm_pu,
	iodc_jtag_ddr_ecc_dq_i,
	iodc_jtag_ddr_ecc_dq_oe_n,
//	iodc_jtag_ddr_ecc_dq_pd,
//	iodc_jtag_ddr_ecc_dq_pu,
	iodc_jtag_ddr_ecc_dqs_i,
	iodc_jtag_ddr_ecc_dqs_oe_n,
//	iodc_jtag_ddr_ecc_dqs_pd,
//	iodc_jtag_ddr_ecc_dqs_pu,
	iodc_jtag_ddr_odt_i,
	iodc_jtag_ddr_odt_oe_n,
//	iodc_jtag_ddr_odt_pd,
//	iodc_jtag_ddr_odt_pu,
	iodc_jtag_ddr_par_i,
	iodc_jtag_ddr_par_oe_n,
//	iodc_jtag_ddr_par_pd,
//	iodc_jtag_ddr_par_pu,
	iodc_jtag_ddr_ras_n_i,
	iodc_jtag_ddr_ras_n_oe_n,
//	iodc_jtag_ddr_ras_n_pd,
//	iodc_jtag_ddr_ras_n_pu,
	iodc_jtag_ddr_reset_n_i,
	iodc_jtag_ddr_reset_n_oe_n,
//	iodc_jtag_ddr_reset_n_pd,
//	iodc_jtag_ddr_reset_n_pu,
	iodc_jtag_ddr_we_n_i,
	iodc_jtag_ddr_we_n_oe_n,
//	iodc_jtag_ddr_we_n_pd,
//	iodc_jtag_ddr_we_n_pu,
//	iodc_jtag_dr3en,
//	iodc_jtag_drvn,
//	iodc_jtag_drvp,
//	iodc_jtag_en,
//	iodc_jtag_gpio_en,
//	iodc_jtag_hv_en,
//	iodc_jtag_odt_ctrl,
//	iodc_jtag_pdm,
//	iodc_jtag_pdn,
//	iodc_jtag_pum,
//	iodc_jtag_smt,
	mc_clk,
	mc_clk_rst_n,
//	phy_scan_clk,
//	phy_scan_en,
//	phy_scan_in_d2f,
//	phy_scan_in_d2r,
//	phy_scan_in_x2f,
//	phy_scan_in_x2r,
//	phy_scan_mode,
//	phy_scan_rst_n,
//	phy_test_iddq,
	r_ddr23phy_reg,
	ddr_addr,
	ddr_bank,
	ddr_cas_n,
	ddr_cke,
	ddr_clk0,
	ddr_clk0_n,
	ddr_cs0_n,
	ddr_dm,
	ddr_dq,
	ddr_dqs,
	ddr_dqs_n,
	ddr_ecc_dm,
	ddr_ecc_dq,
	ddr_ecc_dqs,
	ddr_ecc_dqs_n,
	ddr_odt,
	ddr_ras_n,
	ddr_reset_n,
	ddr_we_n,
	ddr_zq0 
);

output	[31:0]	ahb_hrdata_o;
output		ahb_hready_o;
output	[1:0]	ahb_hresp_o;
output		dram_dfi_ctrlupd_ack;
output	[15:0]	dram_dfi_ecc_rddata_w1;
output	[15:0]	dram_dfi_ecc_rddata_w0;
output		dram_dfi_init_complete;
output	[3:0]	dram_dfi_rddata_valid_w1;
output	[3:0]	dram_dfi_rddata_valid_w0;
output	[63:0]	dram_dfi_rddata_w1;
output	[63:0]	dram_dfi_rddata_w0;
output	[1:0]	dram_dfi_rdlvl_gate_mode;
output	[1:0]	dram_dfi_rdlvl_mode;
output	[39:0]	dram_dfi_rdlvl_resp;
output	[1:0]	dram_dfi_wrlvl_mode;
output	[4:0]	dram_dfi_wrlvl_resp;
output		fp_dfi_ctrlupd_ack;
output		fp_dfi_ecc_rddata_valid_w1;
output		fp_dfi_ecc_rddata_valid_w0;
output	[15:0]	fp_dfi_ecc_rddata_w1;
output	[15:0]	fp_dfi_ecc_rddata_w0;
output		fp_dfi_init_complete;
output	[3:0]	fp_dfi_rddata_valid_w1;
output	[3:0]	fp_dfi_rddata_valid_w0;
output	[63:0]	fp_dfi_rddata_w1;
output	[63:0]	fp_dfi_rddata_w0;
output	[1:0]	fp_dfi_rdlvl_gate_mode;
output	[1:0]	fp_dfi_rdlvl_mode;
output	[39:0]	fp_dfi_rdlvl_resp;
output	[1:0]	fp_dfi_wrlvl_mode;
output	[4:0]	fp_dfi_wrlvl_resp;
output	[15:0]	iodc_jtag_ddr_addr_c;
output	[2:0]	iodc_jtag_ddr_bank_c;
output		iodc_jtag_ddr_cas_n_c;
output		iodc_jtag_ddr_cke_c;
output	[1:0]	iodc_jtag_ddr_clk_c;
output	[1:0]	iodc_jtag_ddr_cs_n_c;
output	[3:0]	iodc_jtag_ddr_dm_c;
output	[31:0]	iodc_jtag_ddr_dq_c;
output	[3:0]	iodc_jtag_ddr_dqs_c;
output		iodc_jtag_ddr_ecc_dm_c;
output	[7:0]	iodc_jtag_ddr_ecc_dq_c;
output		iodc_jtag_ddr_ecc_dqs_c;
output		iodc_jtag_ddr_odt_c;
output		iodc_jtag_ddr_par_c;
output		iodc_jtag_ddr_ras_n_c;
output		iodc_jtag_ddr_reset_n_c;
output		iodc_jtag_ddr_we_n_c;
//output		phy_scan_out_d2f;
//output		phy_scan_out_d2r;
//output		phy_scan_out_x2f;
//output		phy_scan_out_x2r;
output [2047:0]	ro_ddr23phy_reg;
input	[31:0]	ahb_haddr_i;
input	[2:0]	ahb_hburst_i;
input		ahb_hclk;
input		ahb_hready_i;
input		ahb_hresetn;
input		ahb_hsel_i;
input	[2:0]	ahb_hsize_i;
input	[1:0]	ahb_htrans_i;
input	[31:0]	ahb_hwdata_i;
input		ahb_hwrite_i;
input		bypasspll_mc_clk_x4;
//input		dfi_sphy_sel;
input	[19:0]	dram_dfi_addr_p1;
input	[19:0]	dram_dfi_addr_p0;
input	[2:0]	dram_dfi_bank_p1;
input	[2:0]	dram_dfi_bank_p0;
input		dram_dfi_cas_n_p1;
input		dram_dfi_cas_n_p0;
input		dram_dfi_cke_p1;
input		dram_dfi_cke_p0;
input		dram_dfi_cs_n_duplicate_p1;
input		dram_dfi_cs_n_duplicate_p0;
input		dram_dfi_cs_n_p1;
input		dram_dfi_cs_n_p0;
input		dram_dfi_ctrlupd_req;
input		dram_dfi_dram_clk_disable;
input		dram_dfi_ecc_rddata_en_p1;
input		dram_dfi_ecc_rddata_en_p0;
input		dram_dfi_ecc_wrdata_en_p1;
input		dram_dfi_ecc_wrdata_en_p0;
input	[15:0]	dram_dfi_ecc_wrdata_p1;
input	[15:0]	dram_dfi_ecc_wrdata_p0;
input	[1:0]	dram_dfi_ecc_wrmask_p1;
input	[1:0]	dram_dfi_ecc_wrmask_p0;
input		dram_dfi_init_start;
input		dram_dfi_ras_n_p1;
input		dram_dfi_ras_n_p0;
input	[3:0]	dram_dfi_rddata_en_p1;
input	[3:0]	dram_dfi_rddata_en_p0;
input	[15:0]	dram_dfi_rdlvl_delay;
input	[15:0]	dram_dfi_rdlvl_delayn;
input		dram_dfi_rdlvl_edge;
input		dram_dfi_rdlvl_en;
input	[31:0]	dram_dfi_rdlvl_gate_delay;
input		dram_dfi_rdlvl_gate_en;
input		dram_dfi_rdlvl_load;
input		dram_dfi_reset_n_p1;
input		dram_dfi_reset_n_p0;
input		dram_dfi_we_n_p1;
input		dram_dfi_we_n_p0;
input		dram_dfi_wodt_p1;
input		dram_dfi_wodt_p0;
input	[3:0]	dram_dfi_wrdata_en_p1;
input	[3:0]	dram_dfi_wrdata_en_p0;
input	[63:0]	dram_dfi_wrdata_p1;
input	[63:0]	dram_dfi_wrdata_p0;
input	[15:0]	dram_dfi_wrlvl_delay;
input		dram_dfi_wrlvl_en;
input		dram_dfi_wrlvl_load;
input		dram_dfi_wrlvl_strobe;
input	[7:0]	dram_dfi_wrmask_p1;
input	[7:0]	dram_dfi_wrmask_p0;
input	[19:0]	fp_dfi_addr_p1;
input	[19:0]	fp_dfi_addr_p0;
input	[2:0]	fp_dfi_bank_p1;
input	[2:0]	fp_dfi_bank_p0;
input		fp_dfi_cas_n_p1;
input		fp_dfi_cas_n_p0;
input		fp_dfi_cke_p1;
input		fp_dfi_cke_p0;
input		fp_dfi_cs_n_duplicate_p1;
input		fp_dfi_cs_n_duplicate_p0;
input		fp_dfi_cs_n_p1;
input		fp_dfi_cs_n_p0;
input		fp_dfi_ctrlupd_req;
input		fp_dfi_dram_clk_disable;
input		fp_dfi_ecc_rddata_en_p1;
input		fp_dfi_ecc_rddata_en_p0;
input		fp_dfi_ecc_wrdata_en_p1;
input		fp_dfi_ecc_wrdata_en_p0;
input	[15:0]	fp_dfi_ecc_wrdata_p1;
input	[15:0]	fp_dfi_ecc_wrdata_p0;
input	[1:0]	fp_dfi_ecc_wrmask_p1;
input	[1:0]	fp_dfi_ecc_wrmask_p0;
input		fp_dfi_init_start;
input		fp_dfi_ras_n_p1;
input		fp_dfi_ras_n_p0;
input	[3:0]	fp_dfi_rddata_en_p1;
input	[3:0]	fp_dfi_rddata_en_p0;
input	[15:0]	fp_dfi_rdlvl_delay;
input	[15:0]	fp_dfi_rdlvl_delayn;
input		fp_dfi_rdlvl_edge;
input		fp_dfi_rdlvl_en;
input	[31:0]	fp_dfi_rdlvl_gate_delay;
input		fp_dfi_rdlvl_gate_en;
input		fp_dfi_rdlvl_load;
input		fp_dfi_reset_n_p1;
input		fp_dfi_reset_n_p0;
input		fp_dfi_we_n_p1;
input		fp_dfi_we_n_p0;
input		fp_dfi_wodt_p1;
input		fp_dfi_wodt_p0;
input	[3:0]	fp_dfi_wrdata_en_p1;
input	[3:0]	fp_dfi_wrdata_en_p0;
input	[63:0]	fp_dfi_wrdata_p1;
input	[63:0]	fp_dfi_wrdata_p0;
input	[15:0]	fp_dfi_wrlvl_delay;
input		fp_dfi_wrlvl_en;
input		fp_dfi_wrlvl_load;
input		fp_dfi_wrlvl_strobe;
input	[7:0]	fp_dfi_wrmask_p1;
input	[7:0]	fp_dfi_wrmask_p0;
input	[15:0]	iodc_jtag_ddr_addr_i;
input	[15:0]	iodc_jtag_ddr_addr_oe_n;
//input	[15:0]	iodc_jtag_ddr_addr_pd;
//input	[15:0]	iodc_jtag_ddr_addr_pu;
input	[2:0]	iodc_jtag_ddr_bank_i;
input	[2:0]	iodc_jtag_ddr_bank_oe_n;
//input	[2:0]	iodc_jtag_ddr_bank_pd;
//input	[2:0]	iodc_jtag_ddr_bank_pu;
input		iodc_jtag_ddr_cas_n_i;
input		iodc_jtag_ddr_cas_n_oe_n;
//input		iodc_jtag_ddr_cas_n_pd;
//input		iodc_jtag_ddr_cas_n_pu;
input		iodc_jtag_ddr_cke_i;
input		iodc_jtag_ddr_cke_oe_n;
//input		iodc_jtag_ddr_cke_pd;
//input		iodc_jtag_ddr_cke_pu;
input	[1:0]	iodc_jtag_ddr_clk_i;
input	[1:0]	iodc_jtag_ddr_clk_oe_n;
//input	[1:0]	iodc_jtag_ddr_clk_pd;
//input	[1:0]	iodc_jtag_ddr_clk_pu;
input	[1:0]	iodc_jtag_ddr_cs_n_i;
input	[1:0]	iodc_jtag_ddr_cs_n_oe_n;
//input	[1:0]	iodc_jtag_ddr_cs_n_pd;
//input	[1:0]	iodc_jtag_ddr_cs_n_pu;
input	[3:0]	iodc_jtag_ddr_dm_i;
input	[3:0]	iodc_jtag_ddr_dm_oe_n;
//input	[3:0]	iodc_jtag_ddr_dm_pd;
//input	[3:0]	iodc_jtag_ddr_dm_pu;
input	[31:0]	iodc_jtag_ddr_dq_i;
input	[31:0]	iodc_jtag_ddr_dq_oe_n;
//input	[31:0]	iodc_jtag_ddr_dq_pd;
//input	[31:0]	iodc_jtag_ddr_dq_pu;
input	[3:0]	iodc_jtag_ddr_dqs_i;
input	[3:0]	iodc_jtag_ddr_dqs_oe_n;
//input	[3:0]	iodc_jtag_ddr_dqs_pd;
//input	[3:0]	iodc_jtag_ddr_dqs_pu;
input		iodc_jtag_ddr_ecc_dm_i;
input		iodc_jtag_ddr_ecc_dm_oe_n;
//input		iodc_jtag_ddr_ecc_dm_pd;
//input		iodc_jtag_ddr_ecc_dm_pu;
input	[7:0]	iodc_jtag_ddr_ecc_dq_i;
input	[7:0]	iodc_jtag_ddr_ecc_dq_oe_n;
//input	[7:0]	iodc_jtag_ddr_ecc_dq_pd;
//input	[7:0]	iodc_jtag_ddr_ecc_dq_pu;
input		iodc_jtag_ddr_ecc_dqs_i;
input		iodc_jtag_ddr_ecc_dqs_oe_n;
//input		iodc_jtag_ddr_ecc_dqs_pd;
//input		iodc_jtag_ddr_ecc_dqs_pu;
input		iodc_jtag_ddr_odt_i;
input		iodc_jtag_ddr_odt_oe_n;
//input		iodc_jtag_ddr_odt_pd;
//input		iodc_jtag_ddr_odt_pu;
input		iodc_jtag_ddr_par_i;
input		iodc_jtag_ddr_par_oe_n;
//input		iodc_jtag_ddr_par_pd;
//input		iodc_jtag_ddr_par_pu;
input		iodc_jtag_ddr_ras_n_i;
input		iodc_jtag_ddr_ras_n_oe_n;
//input		iodc_jtag_ddr_ras_n_pd;
//input		iodc_jtag_ddr_ras_n_pu;
input		iodc_jtag_ddr_reset_n_i;
input		iodc_jtag_ddr_reset_n_oe_n;
//input		iodc_jtag_ddr_reset_n_pd;
//input		iodc_jtag_ddr_reset_n_pu;
input		iodc_jtag_ddr_we_n_i;
input		iodc_jtag_ddr_we_n_oe_n;
//input		iodc_jtag_ddr_we_n_pd;
//input		iodc_jtag_ddr_we_n_pu;
//input		iodc_jtag_dr3en;
//input	[2:0]	iodc_jtag_drvn;
//input	[2:0]	iodc_jtag_drvp;
//input		iodc_jtag_en;
//input		iodc_jtag_gpio_en;
//input		iodc_jtag_hv_en;
//input	[2:0]	iodc_jtag_odt_ctrl;
//input	[7:0]	iodc_jtag_pdm;
//input		iodc_jtag_pdn;
//input	[7:0]	iodc_jtag_pum;
//input		iodc_jtag_smt;
input		mc_clk;
input		mc_clk_rst_n;
//input		phy_scan_clk;
//input		phy_scan_en;
//input		phy_scan_in_d2f;
//input		phy_scan_in_d2r;
//input		phy_scan_in_x2f;
//input		phy_scan_in_x2r;
//input		phy_scan_mode;
//input		phy_scan_rst_n;
//input		phy_test_iddq;
input [2047:0]	r_ddr23phy_reg;
inout	[15:0]	ddr_addr;
inout	[2:0]	ddr_bank;
inout		ddr_cas_n;
inout		ddr_cke;
inout	[1:0]	ddr_clk0;
inout	[1:0]	ddr_clk0_n;
inout	[1:0]	ddr_cs0_n;
inout	[3:0]	ddr_dm;
inout	[31:0]	ddr_dq;
inout	[3:0]	ddr_dqs;
inout	[3:0]	ddr_dqs_n;
inout		ddr_ecc_dm;
inout	[7:0]	ddr_ecc_dq;
inout		ddr_ecc_dqs;
inout		ddr_ecc_dqs_n;
inout		ddr_odt;
inout		ddr_ras_n;
inout		ddr_reset_n;
inout		ddr_we_n;
inout		ddr_zq0;

parameter phy_test_iddq = 1'b0;
parameter dfi_sphy_sel = 1'b0;
parameter ddr_phy_iso_en = 1'b0;
parameter ddr_phy_pd = 1'b0;

parameter  iodc_jtag_ddr_addr_pd = 16'b0;
parameter  iodc_jtag_ddr_addr_pu = 16'b0;
parameter  iodc_jtag_ddr_bank_pd = 3'b0;
parameter  iodc_jtag_ddr_bank_pu= 3'b0;
parameter  iodc_jtag_ddr_cas_n_pd = 1'b0;
parameter  iodc_jtag_ddr_cas_n_pu = 1'b0;
parameter  iodc_jtag_ddr_cke_pd = 1'b0;
parameter  iodc_jtag_ddr_cke_pu = 1'b0;
parameter  iodc_jtag_ddr_clk_pd = 2'b0;
parameter  iodc_jtag_ddr_clk_pu = 2'b0;
parameter  iodc_jtag_ddr_cs_n_pd = 2'b0;
parameter  iodc_jtag_ddr_cs_n_pu = 2'b0;
parameter  iodc_jtag_ddr_dm_pd = 4'b0;
parameter  iodc_jtag_ddr_dm_pu = 4'b0;
parameter  iodc_jtag_ddr_dq_pd = 32'b0;
parameter  iodc_jtag_ddr_dq_pu = 32'b0;
parameter  iodc_jtag_ddr_dqs_pd = 4'b0;
parameter  iodc_jtag_ddr_dqs_pu = 4'b0;
parameter  iodc_jtag_ddr_ecc_dm_pd = 1'b0;
parameter  iodc_jtag_ddr_ecc_dm_pu = 1'b0;
parameter  iodc_jtag_ddr_ecc_dq_pd = 8'b0;
parameter  iodc_jtag_ddr_ecc_dq_pu = 8'b0;
parameter  iodc_jtag_ddr_ecc_dqs_pd = 1'b0;
parameter  iodc_jtag_ddr_ecc_dqs_pu = 1'b0;
parameter  iodc_jtag_ddr_odt_pd = 1'b0;
parameter  iodc_jtag_ddr_odt_pu = 1'b0;
parameter  iodc_jtag_ddr_par_pd = 1'b0;
parameter  iodc_jtag_ddr_par_pu = 1'b0;
parameter  iodc_jtag_ddr_ras_n_pd = 1'b0;
parameter  iodc_jtag_ddr_ras_n_pu = 1'b0;
parameter  iodc_jtag_ddr_reset_n_pd = 1'b0;
parameter  iodc_jtag_ddr_reset_n_pu = 1'b0;
parameter  iodc_jtag_ddr_we_n_pd = 1'b0;
parameter  iodc_jtag_ddr_we_n_pu = 1'b0;
parameter  iodc_jtag_dr3en = 1'b0;
parameter  iodc_jtag_drvn = 3'b0;
parameter  iodc_jtag_drvp = 3'b0;
parameter  iodc_jtag_en = 1'b0;
parameter  iodc_jtag_gpio_en = 1'b0;
parameter  iodc_jtag_hv_en = 1'b0;
parameter  iodc_jtag_odt_ctrl = 3'b0;
parameter  iodc_jtag_pdm = 8'b0;
parameter  iodc_jtag_pdn = 1'b0;
parameter  iodc_jtag_pum = 8'b0;
parameter  iodc_jtag_smt = 1'b0;

endmodule

// VPERL: GENERATED_END

module SERDES_PHY_V1(
	HP2SP_L3RxCALDetected,
	HP2SP_L3RxGearboxIsSync,
	HP2SP_L3RxOOBCOMINITDet,
	HP2SP_L3RxOOBCOMSASDet,
	HP2SP_L3RxOOBCOMWAKEDet,
	HP2SP_L3RxOOBElecIdle,
	HP2SP_L3RxOvrsmplErr,
	HP2SP_L3RxPIPEPHYStatusRxDet,
	HP2SP_L3RxPIPERxDetected,
	HP2SP_L3RxPRBSErrCnt,
	HP2SP_L3RxPRBSZeroCnt,
	HP2SP_L3RxRecClk,
	HP2SP_L3RxRecClk2,
	HP2SP_L3RxSyncState,
	HP2SP_L3RxUsr8B10BDispErr,
	HP2SP_L3RxUsr8B10BEBCorCnt,
	HP2SP_L3RxUsr8B10BEBStat,
	HP2SP_L3RxUsr8B10BIsComma,
	HP2SP_L3RxUsr8B10BIsK,
	HP2SP_L3RxUsr8B10BNotInTable,
	HP2SP_L3RxUsr8B10BRunDisp,
	HP2SP_L3RxUsr8B10BValid,
	HP2SP_L3RxUsrData,
	HP2SP_L3RxUsrDataValid,
	HP2SP_L3RxUsrGBHeader,
	HP2SP_L3RxUsrGBHeaderValid,
	HP2SP_L3RxUsrGBStartSeq,
	HP2SP_L3TxBufStatus,
	HP2SP_L3TxOutClk,
	HP2SP_L3TxOutClk2,
	HP2SP_L3TxSATAOOBComFinish,
	HP2SP_L3TxUsrGBReady,
	HP2SP_L2RxCALDetected,
	HP2SP_L2RxGearboxIsSync,
	HP2SP_L2RxOOBCOMINITDet,
	HP2SP_L2RxOOBCOMSASDet,
	HP2SP_L2RxOOBCOMWAKEDet,
	HP2SP_L2RxOOBElecIdle,
	HP2SP_L2RxOvrsmplErr,
	HP2SP_L2RxPIPEPHYStatusRxDet,
	HP2SP_L2RxPIPERxDetected,
	HP2SP_L2RxPRBSErrCnt,
	HP2SP_L2RxPRBSZeroCnt,
	HP2SP_L2RxRecClk,
	HP2SP_L2RxRecClk2,
	HP2SP_L2RxSyncState,
	HP2SP_L2RxUsr8B10BDispErr,
	HP2SP_L2RxUsr8B10BEBCorCnt,
	HP2SP_L2RxUsr8B10BEBStat,
	HP2SP_L2RxUsr8B10BIsComma,
	HP2SP_L2RxUsr8B10BIsK,
	HP2SP_L2RxUsr8B10BNotInTable,
	HP2SP_L2RxUsr8B10BRunDisp,
	HP2SP_L2RxUsr8B10BValid,
	HP2SP_L2RxUsrData,
	HP2SP_L2RxUsrDataValid,
	HP2SP_L2RxUsrGBHeader,
	HP2SP_L2RxUsrGBHeaderValid,
	HP2SP_L2RxUsrGBStartSeq,
	HP2SP_L2TxBufStatus,
	HP2SP_L2TxOutClk,
	HP2SP_L2TxOutClk2,
	HP2SP_L2TxSATAOOBComFinish,
	HP2SP_L2TxUsrGBReady,
	HP2SP_L1RxCALDetected,
	HP2SP_L1RxGearboxIsSync,
	HP2SP_L1RxOOBCOMINITDet,
	HP2SP_L1RxOOBCOMSASDet,
	HP2SP_L1RxOOBCOMWAKEDet,
	HP2SP_L1RxOOBElecIdle,
	HP2SP_L1RxOvrsmplErr,
	HP2SP_L1RxPIPEPHYStatusRxDet,
	HP2SP_L1RxPIPERxDetected,
	HP2SP_L1RxPRBSErrCnt,
	HP2SP_L1RxPRBSZeroCnt,
	HP2SP_L1RxRecClk,
	HP2SP_L1RxRecClk2,
	HP2SP_L1RxSyncState,
	HP2SP_L1RxUsr8B10BDispErr,
	HP2SP_L1RxUsr8B10BEBCorCnt,
	HP2SP_L1RxUsr8B10BEBStat,
	HP2SP_L1RxUsr8B10BIsComma,
	HP2SP_L1RxUsr8B10BIsK,
	HP2SP_L1RxUsr8B10BNotInTable,
	HP2SP_L1RxUsr8B10BRunDisp,
	HP2SP_L1RxUsr8B10BValid,
	HP2SP_L1RxUsrData,
	HP2SP_L1RxUsrDataValid,
	HP2SP_L1RxUsrGBHeader,
	HP2SP_L1RxUsrGBHeaderValid,
	HP2SP_L1RxUsrGBStartSeq,
	HP2SP_L1TxBufStatus,
	HP2SP_L1TxOutClk,
	HP2SP_L1TxOutClk2,
	HP2SP_L1TxSATAOOBComFinish,
	HP2SP_L1TxUsrGBReady,
	HP2SP_L0RxCALDetected,
	HP2SP_L0RxGearboxIsSync,
	HP2SP_L0RxOOBCOMINITDet,
	HP2SP_L0RxOOBCOMSASDet,
	HP2SP_L0RxOOBCOMWAKEDet,
	HP2SP_L0RxOOBElecIdle,
	HP2SP_L0RxOvrsmplErr,
	HP2SP_L0RxPIPEPHYStatusRxDet,
	HP2SP_L0RxPIPERxDetected,
	HP2SP_L0RxPRBSErrCnt,
	HP2SP_L0RxPRBSZeroCnt,
	HP2SP_L0RxRecClk,
	HP2SP_L0RxRecClk2,
	HP2SP_L0RxSyncState,
	HP2SP_L0RxUsr8B10BDispErr,
	HP2SP_L0RxUsr8B10BEBCorCnt,
	HP2SP_L0RxUsr8B10BEBStat,
	HP2SP_L0RxUsr8B10BIsComma,
	HP2SP_L0RxUsr8B10BIsK,
	HP2SP_L0RxUsr8B10BNotInTable,
	HP2SP_L0RxUsr8B10BRunDisp,
	HP2SP_L0RxUsr8B10BValid,
	HP2SP_L0RxUsrData,
	HP2SP_L0RxUsrDataValid,
	HP2SP_L0RxUsrGBHeader,
	HP2SP_L0RxUsrGBHeaderValid,
	HP2SP_L0RxUsrGBStartSeq,
	HP2SP_L0TxBufStatus,
	HP2SP_L0TxOutClk,
	HP2SP_L0TxOutClk2,
	HP2SP_L0TxSATAOOBComFinish,
	HP2SP_L0TxUsrGBReady,
	HP2SP_PIPEPhyStatusForce,
	HP2SP_PIPEPhyStatusSoft,
	HP2SP_PowerOnDone,
	HP2SP_RxLDuAlignAcqr,
	HP2SP_SysClk,
	HP2SP_xJTAG_tdo,
	HP2SP_xPLL_DivClk,
	HP2fp_L3RxCALDetected,
	HP2fp_L3RxGearboxIsSync,
	HP2fp_L3RxOOBCOMINITDet,
	HP2fp_L3RxOOBCOMSASDet,
	HP2fp_L3RxOOBCOMWAKEDet,
	HP2fp_L3RxOOBElecIdle,
	HP2fp_L3RxOvrsmplErr,
	HP2fp_L3RxPIPEPHYStatusRxDet,
	HP2fp_L3RxPIPERxDetected,
	HP2fp_L3RxPRBSErrCnt,
	HP2fp_L3RxPRBSZeroCnt,
	HP2fp_L3RxSyncState,
	HP2fp_L3RxUsr8B10BDispErr,
	HP2fp_L3RxUsr8B10BEBCorCnt,
	HP2fp_L3RxUsr8B10BEBStat,
	HP2fp_L3RxUsr8B10BIsComma,
	HP2fp_L3RxUsr8B10BIsK,
	HP2fp_L3RxUsr8B10BNotInTable,
	HP2fp_L3RxUsr8B10BRunDisp,
	HP2fp_L3RxUsr8B10BValid,
	HP2fp_L3RxUsrData,
	HP2fp_L3RxUsrGBHeader,
	HP2fp_L3RxUsrGBHeaderValid,
	HP2fp_L3RxUsrGBStartSeq,
	HP2fp_L3TxBufStatus,
	HP2fp_L3TxSATAOOBComFinish,
	HP2fp_L3TxUsrGBReady,
	HP2fp_L2RxCALDetected,
	HP2fp_L2RxGearboxIsSync,
	HP2fp_L2RxOOBCOMINITDet,
	HP2fp_L2RxOOBCOMSASDet,
	HP2fp_L2RxOOBCOMWAKEDet,
	HP2fp_L2RxOOBElecIdle,
	HP2fp_L2RxOvrsmplErr,
	HP2fp_L2RxPIPEPHYStatusRxDet,
	HP2fp_L2RxPIPERxDetected,
	HP2fp_L2RxPRBSErrCnt,
	HP2fp_L2RxPRBSZeroCnt,
	HP2fp_L2RxSyncState,
	HP2fp_L2RxUsr8B10BDispErr,
	HP2fp_L2RxUsr8B10BEBCorCnt,
	HP2fp_L2RxUsr8B10BEBStat,
	HP2fp_L2RxUsr8B10BIsComma,
	HP2fp_L2RxUsr8B10BIsK,
	HP2fp_L2RxUsr8B10BNotInTable,
	HP2fp_L2RxUsr8B10BRunDisp,
	HP2fp_L2RxUsr8B10BValid,
	HP2fp_L2RxUsrData,
	HP2fp_L2RxUsrGBHeader,
	HP2fp_L2RxUsrGBHeaderValid,
	HP2fp_L2RxUsrGBStartSeq,
	HP2fp_L2TxBufStatus,
	HP2fp_L2TxSATAOOBComFinish,
	HP2fp_L2TxUsrGBReady,
	HP2fp_L1RxCALDetected,
	HP2fp_L1RxGearboxIsSync,
	HP2fp_L1RxOOBCOMINITDet,
	HP2fp_L1RxOOBCOMSASDet,
	HP2fp_L1RxOOBCOMWAKEDet,
	HP2fp_L1RxOOBElecIdle,
	HP2fp_L1RxOvrsmplErr,
	HP2fp_L1RxPIPEPHYStatusRxDet,
	HP2fp_L1RxPIPERxDetected,
	HP2fp_L1RxPRBSErrCnt,
	HP2fp_L1RxPRBSZeroCnt,
	HP2fp_L1RxSyncState,
	HP2fp_L1RxUsr8B10BDispErr,
	HP2fp_L1RxUsr8B10BEBCorCnt,
	HP2fp_L1RxUsr8B10BEBStat,
	HP2fp_L1RxUsr8B10BIsComma,
	HP2fp_L1RxUsr8B10BIsK,
	HP2fp_L1RxUsr8B10BNotInTable,
	HP2fp_L1RxUsr8B10BRunDisp,
	HP2fp_L1RxUsr8B10BValid,
	HP2fp_L1RxUsrData,
	HP2fp_L1RxUsrGBHeader,
	HP2fp_L1RxUsrGBHeaderValid,
	HP2fp_L1RxUsrGBStartSeq,
	HP2fp_L1TxBufStatus,
	HP2fp_L1TxSATAOOBComFinish,
	HP2fp_L1TxUsrGBReady,
	HP2fp_L0RxCALDetected,
	HP2fp_L0RxGearboxIsSync,
	HP2fp_L0RxOOBCOMINITDet,
	HP2fp_L0RxOOBCOMSASDet,
	HP2fp_L0RxOOBCOMWAKEDet,
	HP2fp_L0RxOOBElecIdle,
	HP2fp_L0RxOvrsmplErr,
	HP2fp_L0RxPIPEPHYStatusRxDet,
	HP2fp_L0RxPIPERxDetected,
	HP2fp_L0RxPRBSErrCnt,
	HP2fp_L0RxPRBSZeroCnt,
	HP2fp_L0RxSyncState,
	HP2fp_L0RxUsr8B10BDispErr,
	HP2fp_L0RxUsr8B10BEBCorCnt,
	HP2fp_L0RxUsr8B10BEBStat,
	HP2fp_L0RxUsr8B10BIsComma,
	HP2fp_L0RxUsr8B10BIsK,
	HP2fp_L0RxUsr8B10BNotInTable,
	HP2fp_L0RxUsr8B10BRunDisp,
	HP2fp_L0RxUsr8B10BValid,
	HP2fp_L0RxUsrData,
	HP2fp_L0RxUsrGBHeader,
	HP2fp_L0RxUsrGBHeaderValid,
	HP2fp_L0RxUsrGBStartSeq,
	HP2fp_L0TxBufStatus,
	HP2fp_L0TxSATAOOBComFinish,
	HP2fp_L0TxUsrGBReady,
	HP2fp_PIPEPhyStatusForce,
	HP2fp_PIPEPhyStatusSoft,
	HP2fp_PowerOnDone,
	HP2fp_RxLDuAlignAcqr,
	HP2fp_xPLL_lockdet,
	TSTCK3,
	TSTCK2,
	TSTCK1,
	TSTCK0,
	TXN3,
	TXN2,
	TXN1,
	TXN0,
	TXP3,
	TXP2,
	TXP1,
	TXP0,
	pbus_gnt,
	pbus_rdata,
	REFCLKN,
	REFCLKP,
	RXN3,
	RXN2,
	RXN1,
	RXN0,
	RXP3,
	RXP2,
	RXP1,
	RXP0,
	SP2HP_L3RXClkCorUse,
	SP2HP_L3Rx8B10BDecMComDet,
	SP2HP_L3Rx8B10BDecPComDet,
	SP2HP_L3Rx8B10BUse,
	SP2HP_L3Rx8B10BUserDefCom,
	SP2HP_L3Rx8B10BValidComOnly,
	SP2HP_L3Rx4B5BAlignEn,
	SP2HP_L3Rx4B5BED,
	SP2HP_L3Rx4B5BSD,
	SP2HP_L3Rx4B5BUse,
	SP2HP_L3RxBitReverse,
	SP2HP_L3RxBufClr,
	SP2HP_L3RxBufDepth,
	SP2HP_L3RxBufUse,
	SP2HP_L3RxCAL10BEnable,
	SP2HP_L3RxCALAlignWord,
	SP2HP_L3RxCALDetUse,
	SP2HP_L3RxCALDouble,
	SP2HP_L3RxCALEnMComAlign,
	SP2HP_L3RxCALEnPComAlign,
	SP2HP_L3RxCALMComDet,
	SP2HP_L3RxCALMComValue,
	SP2HP_L3RxCALPComDet,
	SP2HP_L3RxCALPComValue,
	SP2HP_L3RxCALSlide,
	SP2HP_L3RxCALSlideMode,
	SP2HP_L3RxCHBondSeq1,
	SP2HP_L3RxCHBondSeq1En,
	SP2HP_L3RxCHBondSeq1Mask,
	SP2HP_L3RxClkCorAdjLen,
	SP2HP_L3RxClkCorSeq14,
	SP2HP_L3RxClkCorSeq13,
	SP2HP_L3RxClkCorSeq12,
	SP2HP_L3RxClkCorSeq11,
	SP2HP_L3RxClkCorSeq1En,
	SP2HP_L3RxDataWidth,
	SP2HP_L3RxGearboxADJSel,
	SP2HP_L3RxGearboxEnDec,
	SP2HP_L3RxGearboxSlip,
	SP2HP_L3RxGearboxUse,
	SP2HP_L3RxInternalWidth,
	SP2HP_L3RxLDEn,
	SP2HP_L3RxNELClkMuxSel,
	SP2HP_L3RxNLMux,
	SP2HP_L3RxNLMuxWidth,
	SP2HP_L3RxOOBBurstVal,
	SP2HP_L3RxOOBMaxBurst,
	SP2HP_L3RxOOBMaxCOMINIT,
	SP2HP_L3RxOOBMaxCOMSAS,
	SP2HP_L3RxOOBMaxCOMWAKE,
	SP2HP_L3RxOOBMinBurst,
	SP2HP_L3RxOOBMinCOMINIT,
	SP2HP_L3RxOOBMinCOMSAS,
	SP2HP_L3RxOOBMinCOMWAKE,
	SP2HP_L3RxOvrsmplEnAlign,
	SP2HP_L3RxOvrsmplMode,
	SP2HP_L3RxPMux,
	SP2HP_L3RxPRBSCntClr,
	SP2HP_L3RxPRBSTst,
	SP2HP_L3RxPRBSUsr,
	SP2HP_L3RxPRBSWidth,
	SP2HP_L3RxPRBSZCntClr,
	SP2HP_L3RxPolarity,
	SP2HP_L3RxRecClkMuxSel,
	SP2HP_L3RxSyncEn,
	SP2HP_L3RxSyncInvalidIncr,
	SP2HP_L3RxSyncThres,
	SP2HP_L3RxSyncThreshold,
	SP2HP_L3RxUClk2MuxSel,
	SP2HP_L3RxUClkMuxSel,
	SP2HP_L3RxUsrClk,
	SP2HP_L3RxUsrClk2,
	SP2HP_L3Tx8B10BUse,
	SP2HP_L3Tx4B5BUse,
	SP2HP_L3TxBitReverse,
	SP2HP_L3TxBufClr,
	SP2HP_L3TxBufWidth,
	SP2HP_L3TxBufferUse,
	SP2HP_L3TxDMux,
	SP2HP_L3TxDataWidth,
	SP2HP_L3TxElecIdleAdj,
	SP2HP_L3TxFlMux,
	SP2HP_L3TxGearboxFunc,
	SP2HP_L3TxGearboxReadyPre,
	SP2HP_L3TxGearboxUse,
	SP2HP_L3TxInternalWidth,
	SP2HP_L3TxOOBMode,
	SP2HP_L3TxOutClkMuxSel,
	SP2HP_L3TxOvrsmplMode,
	SP2HP_L3TxPCIEBeaconPWidth,
	SP2HP_L3TxPCIEDetectRx,
	SP2HP_L3TxPCIEElecIdle,
	SP2HP_L3TxPClkMuxSel,
	SP2HP_L3TxPMux,
	SP2HP_L3TxPRBSErrCont,
	SP2HP_L3TxPRBSErrOne,
	SP2HP_L3TxPRBSTst,
	SP2HP_L3TxPRBSUsr,
	SP2HP_L3TxPRBSWidth,
	SP2HP_L3TxPolarity,
	SP2HP_L3TxSATAOOBComBurstVal,
	SP2HP_L3TxSATAOOBComRESET,
	SP2HP_L3TxSATAOOBComSAS,
	SP2HP_L3TxSATAOOBComWAKE,
	SP2HP_L3TxSATAOOBType,
	SP2HP_L3TxUClk2MuxSel,
	SP2HP_L3TxUClkMuxSel,
	SP2HP_L3TxUIASmpl,
	SP2HP_L3TxUsr8B10BDataK,
	SP2HP_L3TxUsr8B10BDispMode,
	SP2HP_L3TxUsr8B10BDispVal,
	SP2HP_L3TxUsrClk,
	SP2HP_L3TxUsrClk2,
	SP2HP_L3TxUsrData,
	SP2HP_L3TxUsrGBHeader,
	SP2HP_L3TxUsrGBSequence,
	SP2HP_L3TxUsrGBStartSeq,
	SP2HP_L2RXClkCorUse,
	SP2HP_L2Rx8B10BDecMComDet,
	SP2HP_L2Rx8B10BDecPComDet,
	SP2HP_L2Rx8B10BUse,
	SP2HP_L2Rx8B10BUserDefCom,
	SP2HP_L2Rx8B10BValidComOnly,
	SP2HP_L2Rx4B5BAlignEn,
	SP2HP_L2Rx4B5BED,
	SP2HP_L2Rx4B5BSD,
	SP2HP_L2Rx4B5BUse,
	SP2HP_L2RxBitReverse,
	SP2HP_L2RxBufClr,
	SP2HP_L2RxBufDepth,
	SP2HP_L2RxBufUse,
	SP2HP_L2RxCAL10BEnable,
	SP2HP_L2RxCALAlignWord,
	SP2HP_L2RxCALDetUse,
	SP2HP_L2RxCALDouble,
	SP2HP_L2RxCALEnMComAlign,
	SP2HP_L2RxCALEnPComAlign,
	SP2HP_L2RxCALMComDet,
	SP2HP_L2RxCALMComValue,
	SP2HP_L2RxCALPComDet,
	SP2HP_L2RxCALPComValue,
	SP2HP_L2RxCALSlide,
	SP2HP_L2RxCALSlideMode,
	SP2HP_L2RxCHBondSeq1,
	SP2HP_L2RxCHBondSeq1En,
	SP2HP_L2RxCHBondSeq1Mask,
	SP2HP_L2RxClkCorAdjLen,
	SP2HP_L2RxClkCorSeq14,
	SP2HP_L2RxClkCorSeq13,
	SP2HP_L2RxClkCorSeq12,
	SP2HP_L2RxClkCorSeq11,
	SP2HP_L2RxClkCorSeq1En,
	SP2HP_L2RxDataWidth,
	SP2HP_L2RxGearboxADJSel,
	SP2HP_L2RxGearboxEnDec,
	SP2HP_L2RxGearboxSlip,
	SP2HP_L2RxGearboxUse,
	SP2HP_L2RxInternalWidth,
	SP2HP_L2RxLDEn,
	SP2HP_L2RxNELClkMuxSel,
	SP2HP_L2RxNLMux,
	SP2HP_L2RxNLMuxWidth,
	SP2HP_L2RxOOBBurstVal,
	SP2HP_L2RxOOBMaxBurst,
	SP2HP_L2RxOOBMaxCOMINIT,
	SP2HP_L2RxOOBMaxCOMSAS,
	SP2HP_L2RxOOBMaxCOMWAKE,
	SP2HP_L2RxOOBMinBurst,
	SP2HP_L2RxOOBMinCOMINIT,
	SP2HP_L2RxOOBMinCOMSAS,
	SP2HP_L2RxOOBMinCOMWAKE,
	SP2HP_L2RxOvrsmplEnAlign,
	SP2HP_L2RxOvrsmplMode,
	SP2HP_L2RxPMux,
	SP2HP_L2RxPRBSCntClr,
	SP2HP_L2RxPRBSTst,
	SP2HP_L2RxPRBSUsr,
	SP2HP_L2RxPRBSWidth,
	SP2HP_L2RxPRBSZCntClr,
	SP2HP_L2RxPolarity,
	SP2HP_L2RxRecClkMuxSel,
	SP2HP_L2RxSyncEn,
	SP2HP_L2RxSyncInvalidIncr,
	SP2HP_L2RxSyncThres,
	SP2HP_L2RxSyncThreshold,
	SP2HP_L2RxUClk2MuxSel,
	SP2HP_L2RxUClkMuxSel,
	SP2HP_L2RxUsrClk,
	SP2HP_L2RxUsrClk2,
	SP2HP_L2Tx8B10BUse,
	SP2HP_L2Tx4B5BUse,
	SP2HP_L2TxBitReverse,
	SP2HP_L2TxBufClr,
	SP2HP_L2TxBufWidth,
	SP2HP_L2TxBufferUse,
	SP2HP_L2TxDMux,
	SP2HP_L2TxDataWidth,
	SP2HP_L2TxElecIdleAdj,
	SP2HP_L2TxFlMux,
	SP2HP_L2TxGearboxFunc,
	SP2HP_L2TxGearboxReadyPre,
	SP2HP_L2TxGearboxUse,
	SP2HP_L2TxInternalWidth,
	SP2HP_L2TxOOBMode,
	SP2HP_L2TxOutClkMuxSel,
	SP2HP_L2TxOvrsmplMode,
	SP2HP_L2TxPCIEBeaconPWidth,
	SP2HP_L2TxPCIEDetectRx,
	SP2HP_L2TxPCIEElecIdle,
	SP2HP_L2TxPClkMuxSel,
	SP2HP_L2TxPMux,
	SP2HP_L2TxPRBSErrCont,
	SP2HP_L2TxPRBSErrOne,
	SP2HP_L2TxPRBSTst,
	SP2HP_L2TxPRBSUsr,
	SP2HP_L2TxPRBSWidth,
	SP2HP_L2TxPolarity,
	SP2HP_L2TxSATAOOBComBurstVal,
	SP2HP_L2TxSATAOOBComRESET,
	SP2HP_L2TxSATAOOBComSAS,
	SP2HP_L2TxSATAOOBComWAKE,
	SP2HP_L2TxSATAOOBType,
	SP2HP_L2TxUClk2MuxSel,
	SP2HP_L2TxUClkMuxSel,
	SP2HP_L2TxUIASmpl,
	SP2HP_L2TxUsr8B10BDataK,
	SP2HP_L2TxUsr8B10BDispMode,
	SP2HP_L2TxUsr8B10BDispVal,
	SP2HP_L2TxUsrClk,
	SP2HP_L2TxUsrClk2,
	SP2HP_L2TxUsrData,
	SP2HP_L2TxUsrGBHeader,
	SP2HP_L2TxUsrGBSequence,
	SP2HP_L2TxUsrGBStartSeq,
	SP2HP_L1RXClkCorUse,
	SP2HP_L1Rx8B10BDecMComDet,
	SP2HP_L1Rx8B10BDecPComDet,
	SP2HP_L1Rx8B10BUse,
	SP2HP_L1Rx8B10BUserDefCom,
	SP2HP_L1Rx8B10BValidComOnly,
	SP2HP_L1Rx4B5BAlignEn,
	SP2HP_L1Rx4B5BED,
	SP2HP_L1Rx4B5BSD,
	SP2HP_L1Rx4B5BUse,
	SP2HP_L1RxBitReverse,
	SP2HP_L1RxBufClr,
	SP2HP_L1RxBufDepth,
	SP2HP_L1RxBufUse,
	SP2HP_L1RxCAL10BEnable,
	SP2HP_L1RxCALAlignWord,
	SP2HP_L1RxCALDetUse,
	SP2HP_L1RxCALDouble,
	SP2HP_L1RxCALEnMComAlign,
	SP2HP_L1RxCALEnPComAlign,
	SP2HP_L1RxCALMComDet,
	SP2HP_L1RxCALMComValue,
	SP2HP_L1RxCALPComDet,
	SP2HP_L1RxCALPComValue,
	SP2HP_L1RxCALSlide,
	SP2HP_L1RxCALSlideMode,
	SP2HP_L1RxCHBondSeq1,
	SP2HP_L1RxCHBondSeq1En,
	SP2HP_L1RxCHBondSeq1Mask,
	SP2HP_L1RxClkCorAdjLen,
	SP2HP_L1RxClkCorSeq14,
	SP2HP_L1RxClkCorSeq13,
	SP2HP_L1RxClkCorSeq12,
	SP2HP_L1RxClkCorSeq11,
	SP2HP_L1RxClkCorSeq1En,
	SP2HP_L1RxDataWidth,
	SP2HP_L1RxGearboxADJSel,
	SP2HP_L1RxGearboxEnDec,
	SP2HP_L1RxGearboxSlip,
	SP2HP_L1RxGearboxUse,
	SP2HP_L1RxInternalWidth,
	SP2HP_L1RxLDEn,
	SP2HP_L1RxNELClkMuxSel,
	SP2HP_L1RxNLMux,
	SP2HP_L1RxNLMuxWidth,
	SP2HP_L1RxOOBBurstVal,
	SP2HP_L1RxOOBMaxBurst,
	SP2HP_L1RxOOBMaxCOMINIT,
	SP2HP_L1RxOOBMaxCOMSAS,
	SP2HP_L1RxOOBMaxCOMWAKE,
	SP2HP_L1RxOOBMinBurst,
	SP2HP_L1RxOOBMinCOMINIT,
	SP2HP_L1RxOOBMinCOMSAS,
	SP2HP_L1RxOOBMinCOMWAKE,
	SP2HP_L1RxOvrsmplEnAlign,
	SP2HP_L1RxOvrsmplMode,
	SP2HP_L1RxPMux,
	SP2HP_L1RxPRBSCntClr,
	SP2HP_L1RxPRBSTst,
	SP2HP_L1RxPRBSUsr,
	SP2HP_L1RxPRBSWidth,
	SP2HP_L1RxPRBSZCntClr,
	SP2HP_L1RxPolarity,
	SP2HP_L1RxRecClkMuxSel,
	SP2HP_L1RxSyncEn,
	SP2HP_L1RxSyncInvalidIncr,
	SP2HP_L1RxSyncThres,
	SP2HP_L1RxSyncThreshold,
	SP2HP_L1RxUClk2MuxSel,
	SP2HP_L1RxUClkMuxSel,
	SP2HP_L1RxUsrClk,
	SP2HP_L1RxUsrClk2,
	SP2HP_L1Tx8B10BUse,
	SP2HP_L1Tx4B5BUse,
	SP2HP_L1TxBitReverse,
	SP2HP_L1TxBufClr,
	SP2HP_L1TxBufWidth,
	SP2HP_L1TxBufferUse,
	SP2HP_L1TxDMux,
	SP2HP_L1TxDataWidth,
	SP2HP_L1TxElecIdleAdj,
	SP2HP_L1TxFlMux,
	SP2HP_L1TxGearboxFunc,
	SP2HP_L1TxGearboxReadyPre,
	SP2HP_L1TxGearboxUse,
	SP2HP_L1TxInternalWidth,
	SP2HP_L1TxOOBMode,
	SP2HP_L1TxOutClkMuxSel,
	SP2HP_L1TxOvrsmplMode,
	SP2HP_L1TxPCIEBeaconPWidth,
	SP2HP_L1TxPCIEDetectRx,
	SP2HP_L1TxPCIEElecIdle,
	SP2HP_L1TxPClkMuxSel,
	SP2HP_L1TxPMux,
	SP2HP_L1TxPRBSErrCont,
	SP2HP_L1TxPRBSErrOne,
	SP2HP_L1TxPRBSTst,
	SP2HP_L1TxPRBSUsr,
	SP2HP_L1TxPRBSWidth,
	SP2HP_L1TxPolarity,
	SP2HP_L1TxSATAOOBComBurstVal,
	SP2HP_L1TxSATAOOBComRESET,
	SP2HP_L1TxSATAOOBComSAS,
	SP2HP_L1TxSATAOOBComWAKE,
	SP2HP_L1TxSATAOOBType,
	SP2HP_L1TxUClk2MuxSel,
	SP2HP_L1TxUClkMuxSel,
	SP2HP_L1TxUIASmpl,
	SP2HP_L1TxUsr8B10BDataK,
	SP2HP_L1TxUsr8B10BDispMode,
	SP2HP_L1TxUsr8B10BDispVal,
	SP2HP_L1TxUsrClk,
	SP2HP_L1TxUsrClk2,
	SP2HP_L1TxUsrData,
	SP2HP_L1TxUsrGBHeader,
	SP2HP_L1TxUsrGBSequence,
	SP2HP_L1TxUsrGBStartSeq,
	SP2HP_L0RXClkCorUse,
	SP2HP_L0Rx8B10BDecMComDet,
	SP2HP_L0Rx8B10BDecPComDet,
	SP2HP_L0Rx8B10BUse,
	SP2HP_L0Rx8B10BUserDefCom,
	SP2HP_L0Rx8B10BValidComOnly,
	SP2HP_L0Rx4B5BAlignEn,
	SP2HP_L0Rx4B5BED,
	SP2HP_L0Rx4B5BSD,
	SP2HP_L0Rx4B5BUse,
	SP2HP_L0RxBitReverse,
	SP2HP_L0RxBufClr,
	SP2HP_L0RxBufDepth,
	SP2HP_L0RxBufUse,
	SP2HP_L0RxCAL10BEnable,
	SP2HP_L0RxCALAlignWord,
	SP2HP_L0RxCALDetUse,
	SP2HP_L0RxCALDouble,
	SP2HP_L0RxCALEnMComAlign,
	SP2HP_L0RxCALEnPComAlign,
	SP2HP_L0RxCALMComDet,
	SP2HP_L0RxCALMComValue,
	SP2HP_L0RxCALPComDet,
	SP2HP_L0RxCALPComValue,
	SP2HP_L0RxCALSlide,
	SP2HP_L0RxCALSlideMode,
	SP2HP_L0RxCHBondSeq1,
	SP2HP_L0RxCHBondSeq1En,
	SP2HP_L0RxCHBondSeq1Mask,
	SP2HP_L0RxClkCorAdjLen,
	SP2HP_L0RxClkCorSeq14,
	SP2HP_L0RxClkCorSeq13,
	SP2HP_L0RxClkCorSeq12,
	SP2HP_L0RxClkCorSeq11,
	SP2HP_L0RxClkCorSeq1En,
	SP2HP_L0RxDataWidth,
	SP2HP_L0RxGearboxADJSel,
	SP2HP_L0RxGearboxEnDec,
	SP2HP_L0RxGearboxSlip,
	SP2HP_L0RxGearboxUse,
	SP2HP_L0RxInternalWidth,
	SP2HP_L0RxLDEn,
	SP2HP_L0RxNELClkMuxSel,
	SP2HP_L0RxNLMux,
	SP2HP_L0RxNLMuxWidth,
	SP2HP_L0RxOOBBurstVal,
	SP2HP_L0RxOOBMaxBurst,
	SP2HP_L0RxOOBMaxCOMINIT,
	SP2HP_L0RxOOBMaxCOMSAS,
	SP2HP_L0RxOOBMaxCOMWAKE,
	SP2HP_L0RxOOBMinBurst,
	SP2HP_L0RxOOBMinCOMINIT,
	SP2HP_L0RxOOBMinCOMSAS,
	SP2HP_L0RxOOBMinCOMWAKE,
	SP2HP_L0RxOvrsmplEnAlign,
	SP2HP_L0RxOvrsmplMode,
	SP2HP_L0RxPMux,
	SP2HP_L0RxPRBSCntClr,
	SP2HP_L0RxPRBSTst,
	SP2HP_L0RxPRBSUsr,
	SP2HP_L0RxPRBSWidth,
	SP2HP_L0RxPRBSZCntClr,
	SP2HP_L0RxPolarity,
	SP2HP_L0RxRecClkMuxSel,
	SP2HP_L0RxSyncEn,
	SP2HP_L0RxSyncInvalidIncr,
	SP2HP_L0RxSyncThres,
	SP2HP_L0RxSyncThreshold,
	SP2HP_L0RxUClk2MuxSel,
	SP2HP_L0RxUClkMuxSel,
	SP2HP_L0RxUsrClk,
	SP2HP_L0RxUsrClk2,
	SP2HP_L0Tx8B10BUse,
	SP2HP_L0Tx4B5BUse,
	SP2HP_L0TxBitReverse,
	SP2HP_L0TxBufClr,
	SP2HP_L0TxBufWidth,
	SP2HP_L0TxBufferUse,
	SP2HP_L0TxDMux,
	SP2HP_L0TxDataWidth,
	SP2HP_L0TxElecIdleAdj,
	SP2HP_L0TxFlMux,
	SP2HP_L0TxGearboxFunc,
	SP2HP_L0TxGearboxReadyPre,
	SP2HP_L0TxGearboxUse,
	SP2HP_L0TxInternalWidth,
	SP2HP_L0TxOOBMode,
	SP2HP_L0TxOutClkMuxSel,
	SP2HP_L0TxOvrsmplMode,
	SP2HP_L0TxPCIEBeaconPWidth,
	SP2HP_L0TxPCIEDetectRx,
	SP2HP_L0TxPCIEElecIdle,
	SP2HP_L0TxPClkMuxSel,
	SP2HP_L0TxPMux,
	SP2HP_L0TxPRBSErrCont,
	SP2HP_L0TxPRBSErrOne,
	SP2HP_L0TxPRBSTst,
	SP2HP_L0TxPRBSUsr,
	SP2HP_L0TxPRBSWidth,
	SP2HP_L0TxPolarity,
	SP2HP_L0TxSATAOOBComBurstVal,
	SP2HP_L0TxSATAOOBComRESET,
	SP2HP_L0TxSATAOOBComSAS,
	SP2HP_L0TxSATAOOBComWAKE,
	SP2HP_L0TxSATAOOBType,
	SP2HP_L0TxUClk2MuxSel,
	SP2HP_L0TxUClkMuxSel,
	SP2HP_L0TxUIASmpl,
	SP2HP_L0TxUsr8B10BDataK,
	SP2HP_L0TxUsr8B10BDispMode,
	SP2HP_L0TxUsr8B10BDispVal,
	SP2HP_L0TxUsrClk,
	SP2HP_L0TxUsrClk2,
	SP2HP_L0TxUsrData,
	SP2HP_L0TxUsrGBHeader,
	SP2HP_L0TxUsrGBSequence,
	SP2HP_L0TxUsrGBStartSeq,
	SP2HP_LaneEn,
	SP2HP_PCIEMode,
	SP2HP_PonChgClkT2,
	SP2HP_PonChgClkT1,
	SP2HP_PonDfeCalT,
	SP2HP_PonInitT,
	SP2HP_PonOfstCalHiT,
	SP2HP_PonOfstCalLoT,
	SP2HP_PonPllDetT,
	SP2HP_PonPreDfeCalT,
	SP2HP_PonPrePllDetT,
	SP2HP_PonPreResCalT,
	SP2HP_PonPwrIntvalT,
	SP2HP_PonResCalHiT,
	SP2HP_PonResCalLoT,
	SP2HP_RxUnifClkSel,
	SP2HP_RxX4Mode,
	SP2HP_SSCEnX4,
	SP2HP_SysRstBSel,
	SP2HP_TxDetRxT4,
	SP2HP_TxDetRxT3,
	SP2HP_TxDetRxT2,
	SP2HP_TxDetRxT1,
	SP2HP_TxPhaseAlignT,
	SP2HP_TxX4Mode,
	SP2HP_UsrRst_N,
	SP2HP_UsrRxRst_N,
	SP2HP_UsrTxRst_N,
	SP2HP_xBG_SafeMode,
	SP2HP_xBG_pr200clkmux,
	SP2HP_xBG_pr100BRCal,
	SP2HP_xBG_pr100Rx,
	SP2HP_xBG_pr100Tx,
	SP2HP_xBG_pr100spare,
	SP2HP_xBG_prcal100Rx,
	SP2HP_xBG_prcal100Tx,
	SP2HP_xBG_prcal50Pll,
	SP2HP_xBG_prcal50spare,
	SP2HP_xBG_pwrdnB,
	SP2HP_xBG_trim,
	SP2HP_xCDR3_PIbiasTrim,
	SP2HP_xCDR3_PIcapTrim,
	SP2HP_xCDR3_PdivSelRx,
	SP2HP_xCDR3_SelFourFive,
	SP2HP_xCDR3_clkmode,
	SP2HP_xCDR3_dccen,
	SP2HP_xCDR3_dccfix,
	SP2HP_xCDR3_dcctrim,
	SP2HP_xCDR3_hold,
	SP2HP_xCDR3_inc,
	SP2HP_xCDR3_incF,
	SP2HP_xCDR3_limHF,
	SP2HP_xCDR3_limLF,
	SP2HP_xCDR3_metamode,
	SP2HP_xCDR3_mult2F,
	SP2HP_xCDR3_offs,
	SP2HP_xCDR3_pwrdnB,
	SP2HP_xCDR3_updnsw,
	SP2HP_xCDR2_PIbiasTrim,
	SP2HP_xCDR2_PIcapTrim,
	SP2HP_xCDR2_PdivSelRx,
	SP2HP_xCDR2_SelFourFive,
	SP2HP_xCDR2_clkmode,
	SP2HP_xCDR2_dccen,
	SP2HP_xCDR2_dccfix,
	SP2HP_xCDR2_dcctrim,
	SP2HP_xCDR2_hold,
	SP2HP_xCDR2_inc,
	SP2HP_xCDR2_incF,
	SP2HP_xCDR2_limHF,
	SP2HP_xCDR2_limLF,
	SP2HP_xCDR2_metamode,
	SP2HP_xCDR2_mult2F,
	SP2HP_xCDR2_offs,
	SP2HP_xCDR2_pwrdnB,
	SP2HP_xCDR2_updnsw,
	SP2HP_xCDR1_PIbiasTrim,
	SP2HP_xCDR1_PIcapTrim,
	SP2HP_xCDR1_PdivSelRx,
	SP2HP_xCDR1_SelFourFive,
	SP2HP_xCDR1_clkmode,
	SP2HP_xCDR1_dccen,
	SP2HP_xCDR1_dccfix,
	SP2HP_xCDR1_dcctrim,
	SP2HP_xCDR1_hold,
	SP2HP_xCDR1_inc,
	SP2HP_xCDR1_incF,
	SP2HP_xCDR1_limHF,
	SP2HP_xCDR1_limLF,
	SP2HP_xCDR1_metamode,
	SP2HP_xCDR1_mult2F,
	SP2HP_xCDR1_offs,
	SP2HP_xCDR1_pwrdnB,
	SP2HP_xCDR1_updnsw,
	SP2HP_xCDR0_PIbiasTrim,
	SP2HP_xCDR0_PIcapTrim,
	SP2HP_xCDR0_PdivSelRx,
	SP2HP_xCDR0_SelFourFive,
	SP2HP_xCDR0_clkmode,
	SP2HP_xCDR0_dccen,
	SP2HP_xCDR0_dccfix,
	SP2HP_xCDR0_dcctrim,
	SP2HP_xCDR0_hold,
	SP2HP_xCDR0_inc,
	SP2HP_xCDR0_incF,
	SP2HP_xCDR0_limHF,
	SP2HP_xCDR0_limLF,
	SP2HP_xCDR0_metamode,
	SP2HP_xCDR0_mult2F,
	SP2HP_xCDR0_offs,
	SP2HP_xCDR0_pwrdnB,
	SP2HP_xCDR0_updnsw,
	SP2HP_xCMU_clkmux_pwrdnB,
	SP2HP_xCMU_clkmux_swon,
	SP2HP_xCMU_cur_trim,
	SP2HP_xCMU_pwrdnB,
	SP2HP_xCMU_refclk_sel,
	SP2HP_xCTLE3_Adaps_En,
	SP2HP_xCTLE3_Adaps_inc,
	SP2HP_xCTLE3_memCap,
	SP2HP_xCTLE3_memRes3,
	SP2HP_xCTLE3_memRes2,
	SP2HP_xCTLE3_memRes1,
	SP2HP_xCTLE2_Adaps_En,
	SP2HP_xCTLE2_Adaps_inc,
	SP2HP_xCTLE2_memCap,
	SP2HP_xCTLE2_memRes3,
	SP2HP_xCTLE2_memRes2,
	SP2HP_xCTLE2_memRes1,
	SP2HP_xCTLE1_Adaps_En,
	SP2HP_xCTLE1_Adaps_inc,
	SP2HP_xCTLE1_memCap,
	SP2HP_xCTLE1_memRes3,
	SP2HP_xCTLE1_memRes2,
	SP2HP_xCTLE1_memRes1,
	SP2HP_xCTLE0_Adaps_En,
	SP2HP_xCTLE0_Adaps_inc,
	SP2HP_xCTLE0_memCap,
	SP2HP_xCTLE0_memRes3,
	SP2HP_xCTLE0_memRes2,
	SP2HP_xCTLE0_memRes1,
	SP2HP_xDFE3_Adaps_En,
	SP2HP_xDFE3_AnaClkEn,
	SP2HP_xDFE3_EyeScan_En,
	SP2HP_xDFE3_eqGain,
	SP2HP_xDFE3_isoGain,
	SP2HP_xDFE3_memDly,
	SP2HP_xDFE3_memTap4,
	SP2HP_xDFE3_memTap3,
	SP2HP_xDFE3_memTap2,
	SP2HP_xDFE3_memTap1,
	SP2HP_xDFE3_setDly,
	SP2HP_xDFE3_setEq,
	SP2HP_xDFE3_tapcursel,
	SP2HP_xDFE2_Adaps_En,
	SP2HP_xDFE2_AnaClkEn,
	SP2HP_xDFE2_EyeScan_En,
	SP2HP_xDFE2_eqGain,
	SP2HP_xDFE2_isoGain,
	SP2HP_xDFE2_memDly,
	SP2HP_xDFE2_memTap4,
	SP2HP_xDFE2_memTap3,
	SP2HP_xDFE2_memTap2,
	SP2HP_xDFE2_memTap1,
	SP2HP_xDFE2_setDly,
	SP2HP_xDFE2_setEq,
	SP2HP_xDFE2_tapcursel,
	SP2HP_xDFE1_Adaps_En,
	SP2HP_xDFE1_AnaClkEn,
	SP2HP_xDFE1_EyeScan_En,
	SP2HP_xDFE1_eqGain,
	SP2HP_xDFE1_isoGain,
	SP2HP_xDFE1_memDly,
	SP2HP_xDFE1_memTap4,
	SP2HP_xDFE1_memTap3,
	SP2HP_xDFE1_memTap2,
	SP2HP_xDFE1_memTap1,
	SP2HP_xDFE1_setDly,
	SP2HP_xDFE1_setEq,
	SP2HP_xDFE1_tapcursel,
	SP2HP_xDFE0_Adaps_En,
	SP2HP_xDFE0_AnaClkEn,
	SP2HP_xDFE0_EyeScan_En,
	SP2HP_xDFE0_eqGain,
	SP2HP_xDFE0_isoGain,
	SP2HP_xDFE0_memDly,
	SP2HP_xDFE0_memTap4,
	SP2HP_xDFE0_memTap3,
	SP2HP_xDFE0_memTap2,
	SP2HP_xDFE0_memTap1,
	SP2HP_xDFE0_setDly,
	SP2HP_xDFE0_setEq,
	SP2HP_xDFE0_tapcursel,
	SP2HP_xDFECalEn3_mem,
	SP2HP_xDFECalEn3_sel,
	SP2HP_xDFECalEn2_mem,
	SP2HP_xDFECalEn2_sel,
	SP2HP_xDFECalEn1_mem,
	SP2HP_xDFECalEn1_sel,
	SP2HP_xDFECalEn0_mem,
	SP2HP_xDFECalEn0_sel,
	SP2HP_xJTAG_AC_Signal,
	SP2HP_xJTAG_ClockDR,
	SP2HP_xJTAG_En,
	SP2HP_xJTAG_ShiftDR,
	SP2HP_xJTAG_UpdateDR,
	SP2HP_xJTAG_acmode,
	SP2HP_xJTAG_ini_mem,
	SP2HP_xJTAG_pwrdnB,
	SP2HP_xJTAG_tap_resetB,
	SP2HP_xJTAG_tdi,
	SP2HP_xLane3_farlpbken,
	SP2HP_xLane3_nearlpbken,
	SP2HP_xLane2_farlpbken,
	SP2HP_xLane2_nearlpbken,
	SP2HP_xLane1_farlpbken,
	SP2HP_xLane1_nearlpbken,
	SP2HP_xLane0_farlpbken,
	SP2HP_xLane0_nearlpbken,
	SP2HP_xMisc_pwrdnB,
	SP2HP_xMisc_resetB,
	SP2HP_xOSC_CrntEn,
	SP2HP_xOSC_FSEn,
	SP2HP_xOSC_Rtrim,
	SP2HP_xOSC_pwrdnB,
	SP2HP_xOfstCal3_Ovrd,
	SP2HP_xOfstCal3_inc,
	SP2HP_xOfstCal3_mem,
	SP2HP_xOfstCal3_memCtrl,
	SP2HP_xOfstCal3_memEn,
	SP2HP_xOfstCal3_pwrdnB,
	SP2HP_xOfstCal2_Ovrd,
	SP2HP_xOfstCal2_inc,
	SP2HP_xOfstCal2_mem,
	SP2HP_xOfstCal2_memCtrl,
	SP2HP_xOfstCal2_memEn,
	SP2HP_xOfstCal2_pwrdnB,
	SP2HP_xOfstCal1_Ovrd,
	SP2HP_xOfstCal1_inc,
	SP2HP_xOfstCal1_mem,
	SP2HP_xOfstCal1_memCtrl,
	SP2HP_xOfstCal1_memEn,
	SP2HP_xOfstCal1_pwrdnB,
	SP2HP_xOfstCal0_Ovrd,
	SP2HP_xOfstCal0_inc,
	SP2HP_xOfstCal0_mem,
	SP2HP_xOfstCal0_memCtrl,
	SP2HP_xOfstCal0_memEn,
	SP2HP_xOfstCal0_pwrdnB,
	SP2HP_xPLL_CntlLimit_en,
	SP2HP_xPLL_FBDIV,
	SP2HP_xPLL_LockDet_Force_Lock,
	SP2HP_xPLL_Qpump_2,
	SP2HP_xPLL_Qpump_1,
	SP2HP_xPLL_REFDIV,
	SP2HP_xPLL_VCO_Ctuning,
	SP2HP_xPLL_buf_Itrim,
	SP2HP_xPLL_lockdet_en,
	SP2HP_xPLL_lockdet_period_sel,
	SP2HP_xPLL_lockdet_ppm_sel1,
	SP2HP_xPLL_lockdet_ppm_sel0,
	SP2HP_xPLL_pdivSel,
	SP2HP_xPLL_pwrdnB,
	SP2HP_xPLL_resetB,
	SP2HP_xPLL_selFourFive,
	SP2HP_xRX3_busdivSel,
	SP2HP_xRX3_pwrdnB,
	SP2HP_xRX3_set_phase,
	SP2HP_xRX3_slip_clk,
	SP2HP_xRX3_syncRxToUsrclk,
	SP2HP_xRX3_xrChicoOvrPh5to9,
	SP2HP_xRX3_xrChicoOvrd,
	SP2HP_xRX3_xrChicoOvrdEn,
	SP2HP_xRX2_busdivSel,
	SP2HP_xRX2_pwrdnB,
	SP2HP_xRX2_set_phase,
	SP2HP_xRX2_slip_clk,
	SP2HP_xRX2_syncRxToUsrclk,
	SP2HP_xRX2_xrChicoOvrPh5to9,
	SP2HP_xRX2_xrChicoOvrd,
	SP2HP_xRX2_xrChicoOvrdEn,
	SP2HP_xRX1_busdivSel,
	SP2HP_xRX1_pwrdnB,
	SP2HP_xRX1_set_phase,
	SP2HP_xRX1_slip_clk,
	SP2HP_xRX1_syncRxToUsrclk,
	SP2HP_xRX1_xrChicoOvrPh5to9,
	SP2HP_xRX1_xrChicoOvrd,
	SP2HP_xRX1_xrChicoOvrdEn,
	SP2HP_xRX0_busdivSel,
	SP2HP_xRX0_pwrdnB,
	SP2HP_xRX0_set_phase,
	SP2HP_xRX0_slip_clk,
	SP2HP_xRX0_syncRxToUsrclk,
	SP2HP_xRX0_xrChicoOvrPh5to9,
	SP2HP_xRX0_xrChicoOvrd,
	SP2HP_xRX0_xrChicoOvrdEn,
	SP2HP_xRXAFE3_InCMTrim,
	SP2HP_xRXAFE3_rcvShuntEn,
	SP2HP_xRXAFE3_rcvVssTermEn,
	SP2HP_xRXAFE3_rcvVttTermEn,
	SP2HP_xRXAFE3_termRes50En,
	SP2HP_xRXAFE2_InCMTrim,
	SP2HP_xRXAFE2_rcvShuntEn,
	SP2HP_xRXAFE2_rcvVssTermEn,
	SP2HP_xRXAFE2_rcvVttTermEn,
	SP2HP_xRXAFE2_termRes50En,
	SP2HP_xRXAFE1_InCMTrim,
	SP2HP_xRXAFE1_rcvShuntEn,
	SP2HP_xRXAFE1_rcvVssTermEn,
	SP2HP_xRXAFE1_rcvVttTermEn,
	SP2HP_xRXAFE1_termRes50En,
	SP2HP_xRXAFE0_InCMTrim,
	SP2HP_xRXAFE0_rcvShuntEn,
	SP2HP_xRXAFE0_rcvVssTermEn,
	SP2HP_xRXAFE0_rcvVttTermEn,
	SP2HP_xRXAFE0_termRes50En,
	SP2HP_xRXSquelch3_noSigLevel,
	SP2HP_xRXSquelch3_pwrdnB,
	SP2HP_xRXSquelch2_noSigLevel,
	SP2HP_xRXSquelch2_pwrdnB,
	SP2HP_xRXSquelch1_noSigLevel,
	SP2HP_xRXSquelch1_pwrdnB,
	SP2HP_xRXSquelch0_noSigLevel,
	SP2HP_xRXSquelch0_pwrdnB,
	SP2HP_xResCal_Bg_offset,
	SP2HP_xResCal_LPF_offset,
	SP2HP_xResCal_MemCtrl,
	SP2HP_xResCal_MemEn,
	SP2HP_xResCal_MemRes_Bg,
	SP2HP_xResCal_MemRes_LPF,
	SP2HP_xResCal_MemRes_Rx,
	SP2HP_xResCal_MemRes_Tx,
	SP2HP_xResCal_ResBg_sel,
	SP2HP_xResCal_ResLPF_sel,
	SP2HP_xResCal_ResRx_sel,
	SP2HP_xResCal_ResTx_sel,
	SP2HP_xResCal_Rx_offset,
	SP2HP_xResCal_Tx_offset,
	SP2HP_xTOP_DivOOB,
	SP2HP_xTOP_DivSSC,
	SP2HP_xTOP_DivSYS,
	SP2HP_xTOP_SYSClkSel,
	SP2HP_xTX3_ACCCLK_ROTATEH,
	SP2HP_xTX3_ACC_DIN_SEL,
	SP2HP_xTX3_ACC_NSEL,
	SP2HP_xTX3_ACC_OVERRIDE,
	SP2HP_xTX3_ACC_OVERRIDE_EN,
	SP2HP_xTX3_ACC_ROTATE,
	SP2HP_xTX3_ACC_UPDNSW,
	SP2HP_xTX3_Clk_pwrdnB,
	SP2HP_xTX3_DrvPostCursor,
	SP2HP_xTX3_DrvPreCursor,
	SP2HP_xTX3_Drv_pwrdnB,
	SP2HP_xTX3_Drvbiastrim,
	SP2HP_xTX3_Drvswing,
	SP2HP_xTX3_PI_captrim,
	SP2HP_xTX3_PI_pwrdnB,
	SP2HP_xTX3_PIbiasTrim,
	SP2HP_xTX3_Resl_En,
	SP2HP_xTX3_SSC_EN,
	SP2HP_xTX3_SSC_OVERRIDE,
	SP2HP_xTX3_SSC_OVERRIDE_EN,
	SP2HP_xTX3_SSC_TSEL,
	SP2HP_xTX3_Ser_pwrdnB,
	SP2HP_xTX3_Serbiastrim,
	SP2HP_xTX3_Vreftrim,
	SP2HP_xTX3_activepkEn,
	SP2HP_xTX3_busdivSel,
	SP2HP_xTX3_chico_cksel,
	SP2HP_xTX3_chico_pwrdnB,
	SP2HP_xTX3_ctune,
	SP2HP_xTX3_dccbiastrim,
	SP2HP_xTX3_dccerrtrim,
	SP2HP_xTX3_dccfix,
	SP2HP_xTX3_gmtune,
	SP2HP_xTX3_ovsdivEn,
	SP2HP_xTX3_pdivSel,
	SP2HP_xTX3_pwrdnB,
	SP2HP_xTX3_selFourFive,
	SP2HP_xTX3_sendidle,
	SP2HP_xTX3_syncTxToUsrclk,
	SP2HP_xTX3_tdccEn,
	SP2HP_xTX3_tdccovrd,
	SP2HP_xTX2_ACCCLK_ROTATEH,
	SP2HP_xTX2_ACC_DIN_SEL,
	SP2HP_xTX2_ACC_NSEL,
	SP2HP_xTX2_ACC_OVERRIDE,
	SP2HP_xTX2_ACC_OVERRIDE_EN,
	SP2HP_xTX2_ACC_ROTATE,
	SP2HP_xTX2_ACC_UPDNSW,
	SP2HP_xTX2_Clk_pwrdnB,
	SP2HP_xTX2_DrvPostCursor,
	SP2HP_xTX2_DrvPreCursor,
	SP2HP_xTX2_Drv_pwrdnB,
	SP2HP_xTX2_Drvbiastrim,
	SP2HP_xTX2_Drvswing,
	SP2HP_xTX2_PI_captrim,
	SP2HP_xTX2_PI_pwrdnB,
	SP2HP_xTX2_PIbiasTrim,
	SP2HP_xTX2_Resl_En,
	SP2HP_xTX2_SSC_EN,
	SP2HP_xTX2_SSC_OVERRIDE,
	SP2HP_xTX2_SSC_OVERRIDE_EN,
	SP2HP_xTX2_SSC_TSEL,
	SP2HP_xTX2_Ser_pwrdnB,
	SP2HP_xTX2_Serbiastrim,
	SP2HP_xTX2_Vreftrim,
	SP2HP_xTX2_activepkEn,
	SP2HP_xTX2_busdivSel,
	SP2HP_xTX2_chico_cksel,
	SP2HP_xTX2_chico_pwrdnB,
	SP2HP_xTX2_ctune,
	SP2HP_xTX2_dccbiastrim,
	SP2HP_xTX2_dccerrtrim,
	SP2HP_xTX2_dccfix,
	SP2HP_xTX2_gmtune,
	SP2HP_xTX2_ovsdivEn,
	SP2HP_xTX2_pdivSel,
	SP2HP_xTX2_pwrdnB,
	SP2HP_xTX2_selFourFive,
	SP2HP_xTX2_sendidle,
	SP2HP_xTX2_syncTxToUsrclk,
	SP2HP_xTX2_tdccEn,
	SP2HP_xTX2_tdccovrd,
	SP2HP_xTX1_ACCCLK_ROTATEH,
	SP2HP_xTX1_ACC_DIN_SEL,
	SP2HP_xTX1_ACC_NSEL,
	SP2HP_xTX1_ACC_OVERRIDE,
	SP2HP_xTX1_ACC_OVERRIDE_EN,
	SP2HP_xTX1_ACC_ROTATE,
	SP2HP_xTX1_ACC_UPDNSW,
	SP2HP_xTX1_Clk_pwrdnB,
	SP2HP_xTX1_DrvPostCursor,
	SP2HP_xTX1_DrvPreCursor,
	SP2HP_xTX1_Drv_pwrdnB,
	SP2HP_xTX1_Drvbiastrim,
	SP2HP_xTX1_Drvswing,
	SP2HP_xTX1_PI_captrim,
	SP2HP_xTX1_PI_pwrdnB,
	SP2HP_xTX1_PIbiasTrim,
	SP2HP_xTX1_Resl_En,
	SP2HP_xTX1_SSC_EN,
	SP2HP_xTX1_SSC_OVERRIDE,
	SP2HP_xTX1_SSC_OVERRIDE_EN,
	SP2HP_xTX1_SSC_TSEL,
	SP2HP_xTX1_Ser_pwrdnB,
	SP2HP_xTX1_Serbiastrim,
	SP2HP_xTX1_Vreftrim,
	SP2HP_xTX1_activepkEn,
	SP2HP_xTX1_busdivSel,
	SP2HP_xTX1_chico_cksel,
	SP2HP_xTX1_chico_pwrdnB,
	SP2HP_xTX1_ctune,
	SP2HP_xTX1_dccbiastrim,
	SP2HP_xTX1_dccerrtrim,
	SP2HP_xTX1_dccfix,
	SP2HP_xTX1_gmtune,
	SP2HP_xTX1_ovsdivEn,
	SP2HP_xTX1_pdivSel,
	SP2HP_xTX1_pwrdnB,
	SP2HP_xTX1_selFourFive,
	SP2HP_xTX1_sendidle,
	SP2HP_xTX1_syncTxToUsrclk,
	SP2HP_xTX1_tdccEn,
	SP2HP_xTX1_tdccovrd,
	SP2HP_xTX0_ACCCLK_ROTATEH,
	SP2HP_xTX0_ACC_DIN_SEL,
	SP2HP_xTX0_ACC_NSEL,
	SP2HP_xTX0_ACC_OVERRIDE,
	SP2HP_xTX0_ACC_OVERRIDE_EN,
	SP2HP_xTX0_ACC_ROTATE,
	SP2HP_xTX0_ACC_UPDNSW,
	SP2HP_xTX0_Clk_pwrdnB,
	SP2HP_xTX0_DrvPostCursor,
	SP2HP_xTX0_DrvPreCursor,
	SP2HP_xTX0_Drv_pwrdnB,
	SP2HP_xTX0_Drvbiastrim,
	SP2HP_xTX0_Drvswing,
	SP2HP_xTX0_PI_captrim,
	SP2HP_xTX0_PI_pwrdnB,
	SP2HP_xTX0_PIbiasTrim,
	SP2HP_xTX0_Resl_En,
	SP2HP_xTX0_SSC_EN,
	SP2HP_xTX0_SSC_OVERRIDE,
	SP2HP_xTX0_SSC_OVERRIDE_EN,
	SP2HP_xTX0_SSC_TSEL,
	SP2HP_xTX0_Ser_pwrdnB,
	SP2HP_xTX0_Serbiastrim,
	SP2HP_xTX0_Vreftrim,
	SP2HP_xTX0_activepkEn,
	SP2HP_xTX0_busdivSel,
	SP2HP_xTX0_chico_cksel,
	SP2HP_xTX0_chico_pwrdnB,
	SP2HP_xTX0_ctune,
	SP2HP_xTX0_dccbiastrim,
	SP2HP_xTX0_dccerrtrim,
	SP2HP_xTX0_dccfix,
	SP2HP_xTX0_gmtune,
	SP2HP_xTX0_ovsdivEn,
	SP2HP_xTX0_pdivSel,
	SP2HP_xTX0_pwrdnB,
	SP2HP_xTX0_selFourFive,
	SP2HP_xTX0_sendidle,
	SP2HP_xTX0_syncTxToUsrclk,
	SP2HP_xTX0_tdccEn,
	SP2HP_xTX0_tdccovrd,
	SP2HP_xTX_SSC_Align,
	clk_p,
	fp2HP_L3RxBufClr,
	fp2HP_L3RxCALSlide,
	fp2HP_L3RxGearboxSlip,
	fp2HP_L3RxPRBSCntClr,
	fp2HP_L3RxPRBSTst,
	fp2HP_L3RxPRBSZCntClr,
	fp2HP_L3RxPolarity,
	fp2HP_L3TxBitReverse,
	fp2HP_L3TxBufClr,
	fp2HP_L3TxDMux,
	fp2HP_L3TxElecIdleAdj,
	fp2HP_L3TxFlMux,
	fp2HP_L3TxPCIEDetectRx,
	fp2HP_L3TxPCIEElecIdle,
	fp2HP_L3TxPMux,
	fp2HP_L3TxPRBSErrCont,
	fp2HP_L3TxPRBSErrOne,
	fp2HP_L3TxPRBSTst,
	fp2HP_L3TxPolarity,
	fp2HP_L3TxSATAOOBComRESET,
	fp2HP_L3TxSATAOOBComSAS,
	fp2HP_L3TxSATAOOBComWAKE,
	fp2HP_L3TxUsr8B10BDataK,
	fp2HP_L3TxUsr8B10BDispMode,
	fp2HP_L3TxUsr8B10BDispVal,
	fp2HP_L3TxUsrData,
	fp2HP_L3TxUsrGBHeader,
	fp2HP_L3TxUsrGBSequence,
	fp2HP_L3TxUsrGBStartSeq,
	fp2HP_L2RxBufClr,
	fp2HP_L2RxCALSlide,
	fp2HP_L2RxGearboxSlip,
	fp2HP_L2RxPRBSCntClr,
	fp2HP_L2RxPRBSTst,
	fp2HP_L2RxPRBSZCntClr,
	fp2HP_L2RxPolarity,
	fp2HP_L2TxBitReverse,
	fp2HP_L2TxBufClr,
	fp2HP_L2TxDMux,
	fp2HP_L2TxElecIdleAdj,
	fp2HP_L2TxFlMux,
	fp2HP_L2TxPCIEDetectRx,
	fp2HP_L2TxPCIEElecIdle,
	fp2HP_L2TxPMux,
	fp2HP_L2TxPRBSErrCont,
	fp2HP_L2TxPRBSErrOne,
	fp2HP_L2TxPRBSTst,
	fp2HP_L2TxPolarity,
	fp2HP_L2TxSATAOOBComRESET,
	fp2HP_L2TxSATAOOBComSAS,
	fp2HP_L2TxSATAOOBComWAKE,
	fp2HP_L2TxUsr8B10BDataK,
	fp2HP_L2TxUsr8B10BDispMode,
	fp2HP_L2TxUsr8B10BDispVal,
	fp2HP_L2TxUsrData,
	fp2HP_L2TxUsrGBHeader,
	fp2HP_L2TxUsrGBSequence,
	fp2HP_L2TxUsrGBStartSeq,
	fp2HP_L1RxBufClr,
	fp2HP_L1RxCALSlide,
	fp2HP_L1RxGearboxSlip,
	fp2HP_L1RxPRBSCntClr,
	fp2HP_L1RxPRBSTst,
	fp2HP_L1RxPRBSZCntClr,
	fp2HP_L1RxPolarity,
	fp2HP_L1TxBitReverse,
	fp2HP_L1TxBufClr,
	fp2HP_L1TxDMux,
	fp2HP_L1TxElecIdleAdj,
	fp2HP_L1TxFlMux,
	fp2HP_L1TxPCIEDetectRx,
	fp2HP_L1TxPCIEElecIdle,
	fp2HP_L1TxPMux,
	fp2HP_L1TxPRBSErrCont,
	fp2HP_L1TxPRBSErrOne,
	fp2HP_L1TxPRBSTst,
	fp2HP_L1TxPolarity,
	fp2HP_L1TxSATAOOBComRESET,
	fp2HP_L1TxSATAOOBComSAS,
	fp2HP_L1TxSATAOOBComWAKE,
	fp2HP_L1TxUsr8B10BDataK,
	fp2HP_L1TxUsr8B10BDispMode,
	fp2HP_L1TxUsr8B10BDispVal,
	fp2HP_L1TxUsrData,
	fp2HP_L1TxUsrGBHeader,
	fp2HP_L1TxUsrGBSequence,
	fp2HP_L1TxUsrGBStartSeq,
	fp2HP_L0RxBufClr,
	fp2HP_L0RxCALSlide,
	fp2HP_L0RxGearboxSlip,
	fp2HP_L0RxPRBSCntClr,
	fp2HP_L0RxPRBSTst,
	fp2HP_L0RxPRBSZCntClr,
	fp2HP_L0RxPolarity,
	fp2HP_L0TxBitReverse,
	fp2HP_L0TxBufClr,
	fp2HP_L0TxDMux,
	fp2HP_L0TxElecIdleAdj,
	fp2HP_L0TxFlMux,
	fp2HP_L0TxPCIEDetectRx,
	fp2HP_L0TxPCIEElecIdle,
	fp2HP_L0TxPMux,
	fp2HP_L0TxPRBSErrCont,
	fp2HP_L0TxPRBSErrOne,
	fp2HP_L0TxPRBSTst,
	fp2HP_L0TxPolarity,
	fp2HP_L0TxSATAOOBComRESET,
	fp2HP_L0TxSATAOOBComSAS,
	fp2HP_L0TxSATAOOBComWAKE,
	fp2HP_L0TxUsr8B10BDataK,
	fp2HP_L0TxUsr8B10BDispMode,
	fp2HP_L0TxUsr8B10BDispVal,
	fp2HP_L0TxUsrData,
	fp2HP_L0TxUsrGBHeader,
	fp2HP_L0TxUsrGBSequence,
	fp2HP_L0TxUsrGBStartSeq,
	fp2HP_UsrRst_N,
	fp2HP_UsrRxRst_N,
	fp2HP_UsrTxRst_N,
	fp2HP_pcs_usr_resetB,
	pbus_addr,
	pbus_req,
	pbus_wdata,
	pbus_write,
	rst_p_n,
	xCMU_grefclk
);

output		HP2SP_L3RxCALDetected;
output		HP2SP_L3RxGearboxIsSync;
output		HP2SP_L3RxOOBCOMINITDet;
output		HP2SP_L3RxOOBCOMSASDet;
output		HP2SP_L3RxOOBCOMWAKEDet;
output		HP2SP_L3RxOOBElecIdle;
output		HP2SP_L3RxOvrsmplErr;
output		HP2SP_L3RxPIPEPHYStatusRxDet;
output		HP2SP_L3RxPIPERxDetected;
output	[15:0]	HP2SP_L3RxPRBSErrCnt;
output	[15:0]	HP2SP_L3RxPRBSZeroCnt;
output		HP2SP_L3RxRecClk;
output		HP2SP_L3RxRecClk2;
output	[1:0]	HP2SP_L3RxSyncState;
output	[7:0]	HP2SP_L3RxUsr8B10BDispErr;
output	[11:0]	HP2SP_L3RxUsr8B10BEBCorCnt;
output	[11:0]	HP2SP_L3RxUsr8B10BEBStat;
output	[7:0]	HP2SP_L3RxUsr8B10BIsComma;
output	[7:0]	HP2SP_L3RxUsr8B10BIsK;
output	[7:0]	HP2SP_L3RxUsr8B10BNotInTable;
output	[7:0]	HP2SP_L3RxUsr8B10BRunDisp;
output		HP2SP_L3RxUsr8B10BValid;
output	[79:0]	HP2SP_L3RxUsrData;
output		HP2SP_L3RxUsrDataValid;
output	[2:0]	HP2SP_L3RxUsrGBHeader;
output		HP2SP_L3RxUsrGBHeaderValid;
output		HP2SP_L3RxUsrGBStartSeq;
output	[2:0]	HP2SP_L3TxBufStatus;
output		HP2SP_L3TxOutClk;
output		HP2SP_L3TxOutClk2;
output		HP2SP_L3TxSATAOOBComFinish;
output		HP2SP_L3TxUsrGBReady;
output		HP2SP_L2RxCALDetected;
output		HP2SP_L2RxGearboxIsSync;
output		HP2SP_L2RxOOBCOMINITDet;
output		HP2SP_L2RxOOBCOMSASDet;
output		HP2SP_L2RxOOBCOMWAKEDet;
output		HP2SP_L2RxOOBElecIdle;
output		HP2SP_L2RxOvrsmplErr;
output		HP2SP_L2RxPIPEPHYStatusRxDet;
output		HP2SP_L2RxPIPERxDetected;
output	[15:0]	HP2SP_L2RxPRBSErrCnt;
output	[15:0]	HP2SP_L2RxPRBSZeroCnt;
output		HP2SP_L2RxRecClk;
output		HP2SP_L2RxRecClk2;
output	[1:0]	HP2SP_L2RxSyncState;
output	[7:0]	HP2SP_L2RxUsr8B10BDispErr;
output	[11:0]	HP2SP_L2RxUsr8B10BEBCorCnt;
output	[11:0]	HP2SP_L2RxUsr8B10BEBStat;
output	[7:0]	HP2SP_L2RxUsr8B10BIsComma;
output	[7:0]	HP2SP_L2RxUsr8B10BIsK;
output	[7:0]	HP2SP_L2RxUsr8B10BNotInTable;
output	[7:0]	HP2SP_L2RxUsr8B10BRunDisp;
output		HP2SP_L2RxUsr8B10BValid;
output	[79:0]	HP2SP_L2RxUsrData;
output		HP2SP_L2RxUsrDataValid;
output	[2:0]	HP2SP_L2RxUsrGBHeader;
output		HP2SP_L2RxUsrGBHeaderValid;
output		HP2SP_L2RxUsrGBStartSeq;
output	[2:0]	HP2SP_L2TxBufStatus;
output		HP2SP_L2TxOutClk;
output		HP2SP_L2TxOutClk2;
output		HP2SP_L2TxSATAOOBComFinish;
output		HP2SP_L2TxUsrGBReady;
output		HP2SP_L1RxCALDetected;
output		HP2SP_L1RxGearboxIsSync;
output		HP2SP_L1RxOOBCOMINITDet;
output		HP2SP_L1RxOOBCOMSASDet;
output		HP2SP_L1RxOOBCOMWAKEDet;
output		HP2SP_L1RxOOBElecIdle;
output		HP2SP_L1RxOvrsmplErr;
output		HP2SP_L1RxPIPEPHYStatusRxDet;
output		HP2SP_L1RxPIPERxDetected;
output	[15:0]	HP2SP_L1RxPRBSErrCnt;
output	[15:0]	HP2SP_L1RxPRBSZeroCnt;
output		HP2SP_L1RxRecClk;
output		HP2SP_L1RxRecClk2;
output	[1:0]	HP2SP_L1RxSyncState;
output	[7:0]	HP2SP_L1RxUsr8B10BDispErr;
output	[11:0]	HP2SP_L1RxUsr8B10BEBCorCnt;
output	[11:0]	HP2SP_L1RxUsr8B10BEBStat;
output	[7:0]	HP2SP_L1RxUsr8B10BIsComma;
output	[7:0]	HP2SP_L1RxUsr8B10BIsK;
output	[7:0]	HP2SP_L1RxUsr8B10BNotInTable;
output	[7:0]	HP2SP_L1RxUsr8B10BRunDisp;
output		HP2SP_L1RxUsr8B10BValid;
output	[79:0]	HP2SP_L1RxUsrData;
output		HP2SP_L1RxUsrDataValid;
output	[2:0]	HP2SP_L1RxUsrGBHeader;
output		HP2SP_L1RxUsrGBHeaderValid;
output		HP2SP_L1RxUsrGBStartSeq;
output	[2:0]	HP2SP_L1TxBufStatus;
output		HP2SP_L1TxOutClk;
output		HP2SP_L1TxOutClk2;
output		HP2SP_L1TxSATAOOBComFinish;
output		HP2SP_L1TxUsrGBReady;
output		HP2SP_L0RxCALDetected;
output		HP2SP_L0RxGearboxIsSync;
output		HP2SP_L0RxOOBCOMINITDet;
output		HP2SP_L0RxOOBCOMSASDet;
output		HP2SP_L0RxOOBCOMWAKEDet;
output		HP2SP_L0RxOOBElecIdle;
output		HP2SP_L0RxOvrsmplErr;
output		HP2SP_L0RxPIPEPHYStatusRxDet;
output		HP2SP_L0RxPIPERxDetected;
output	[15:0]	HP2SP_L0RxPRBSErrCnt;
output	[15:0]	HP2SP_L0RxPRBSZeroCnt;
output		HP2SP_L0RxRecClk;
output		HP2SP_L0RxRecClk2;
output	[1:0]	HP2SP_L0RxSyncState;
output	[7:0]	HP2SP_L0RxUsr8B10BDispErr;
output	[11:0]	HP2SP_L0RxUsr8B10BEBCorCnt;
output	[11:0]	HP2SP_L0RxUsr8B10BEBStat;
output	[7:0]	HP2SP_L0RxUsr8B10BIsComma;
output	[7:0]	HP2SP_L0RxUsr8B10BIsK;
output	[7:0]	HP2SP_L0RxUsr8B10BNotInTable;
output	[7:0]	HP2SP_L0RxUsr8B10BRunDisp;
output		HP2SP_L0RxUsr8B10BValid;
output	[79:0]	HP2SP_L0RxUsrData;
output		HP2SP_L0RxUsrDataValid;
output	[2:0]	HP2SP_L0RxUsrGBHeader;
output		HP2SP_L0RxUsrGBHeaderValid;
output		HP2SP_L0RxUsrGBStartSeq;
output	[2:0]	HP2SP_L0TxBufStatus;
output		HP2SP_L0TxOutClk;
output		HP2SP_L0TxOutClk2;
output		HP2SP_L0TxSATAOOBComFinish;
output		HP2SP_L0TxUsrGBReady;
output		HP2SP_PIPEPhyStatusForce;
output		HP2SP_PIPEPhyStatusSoft;
output		HP2SP_PowerOnDone;
output		HP2SP_RxLDuAlignAcqr;
output		HP2SP_SysClk;
output		HP2SP_xJTAG_tdo;
output		HP2SP_xPLL_DivClk;
output	[0:0]	HP2fp_L3RxCALDetected;
output	[0:0]	HP2fp_L3RxGearboxIsSync;
output	[0:0]	HP2fp_L3RxOOBCOMINITDet;
output	[0:0]	HP2fp_L3RxOOBCOMSASDet;
output	[0:0]	HP2fp_L3RxOOBCOMWAKEDet;
output	[0:0]	HP2fp_L3RxOOBElecIdle;
output	[0:0]	HP2fp_L3RxOvrsmplErr;
output	[0:0]	HP2fp_L3RxPIPEPHYStatusRxDet;
output	[0:0]	HP2fp_L3RxPIPERxDetected;
output	[15:0]	HP2fp_L3RxPRBSErrCnt;
output	[15:0]	HP2fp_L3RxPRBSZeroCnt;
output	[1:0]	HP2fp_L3RxSyncState;
output	[7:0]	HP2fp_L3RxUsr8B10BDispErr;
output	[11:0]	HP2fp_L3RxUsr8B10BEBCorCnt;
output	[11:0]	HP2fp_L3RxUsr8B10BEBStat;
output	[7:0]	HP2fp_L3RxUsr8B10BIsComma;
output	[7:0]	HP2fp_L3RxUsr8B10BIsK;
output	[7:0]	HP2fp_L3RxUsr8B10BNotInTable;
output	[7:0]	HP2fp_L3RxUsr8B10BRunDisp;
output	[0:0]	HP2fp_L3RxUsr8B10BValid;
output	[79:0]	HP2fp_L3RxUsrData;
output	[2:0]	HP2fp_L3RxUsrGBHeader;
output	[0:0]	HP2fp_L3RxUsrGBHeaderValid;
output	[0:0]	HP2fp_L3RxUsrGBStartSeq;
output	[2:0]	HP2fp_L3TxBufStatus;
output	[0:0]	HP2fp_L3TxSATAOOBComFinish;
output	[0:0]	HP2fp_L3TxUsrGBReady;
output	[0:0]	HP2fp_L2RxCALDetected;
output	[0:0]	HP2fp_L2RxGearboxIsSync;
output	[0:0]	HP2fp_L2RxOOBCOMINITDet;
output	[0:0]	HP2fp_L2RxOOBCOMSASDet;
output	[0:0]	HP2fp_L2RxOOBCOMWAKEDet;
output	[0:0]	HP2fp_L2RxOOBElecIdle;
output	[0:0]	HP2fp_L2RxOvrsmplErr;
output	[0:0]	HP2fp_L2RxPIPEPHYStatusRxDet;
output	[0:0]	HP2fp_L2RxPIPERxDetected;
output	[15:0]	HP2fp_L2RxPRBSErrCnt;
output	[15:0]	HP2fp_L2RxPRBSZeroCnt;
output	[1:0]	HP2fp_L2RxSyncState;
output	[7:0]	HP2fp_L2RxUsr8B10BDispErr;
output	[11:0]	HP2fp_L2RxUsr8B10BEBCorCnt;
output	[11:0]	HP2fp_L2RxUsr8B10BEBStat;
output	[7:0]	HP2fp_L2RxUsr8B10BIsComma;
output	[7:0]	HP2fp_L2RxUsr8B10BIsK;
output	[7:0]	HP2fp_L2RxUsr8B10BNotInTable;
output	[7:0]	HP2fp_L2RxUsr8B10BRunDisp;
output	[0:0]	HP2fp_L2RxUsr8B10BValid;
output	[79:0]	HP2fp_L2RxUsrData;
output	[2:0]	HP2fp_L2RxUsrGBHeader;
output	[0:0]	HP2fp_L2RxUsrGBHeaderValid;
output	[0:0]	HP2fp_L2RxUsrGBStartSeq;
output	[2:0]	HP2fp_L2TxBufStatus;
output	[0:0]	HP2fp_L2TxSATAOOBComFinish;
output	[0:0]	HP2fp_L2TxUsrGBReady;
output	[0:0]	HP2fp_L1RxCALDetected;
output	[0:0]	HP2fp_L1RxGearboxIsSync;
output	[0:0]	HP2fp_L1RxOOBCOMINITDet;
output	[0:0]	HP2fp_L1RxOOBCOMSASDet;
output	[0:0]	HP2fp_L1RxOOBCOMWAKEDet;
output	[0:0]	HP2fp_L1RxOOBElecIdle;
output	[0:0]	HP2fp_L1RxOvrsmplErr;
output	[0:0]	HP2fp_L1RxPIPEPHYStatusRxDet;
output	[0:0]	HP2fp_L1RxPIPERxDetected;
output	[15:0]	HP2fp_L1RxPRBSErrCnt;
output	[15:0]	HP2fp_L1RxPRBSZeroCnt;
output	[1:0]	HP2fp_L1RxSyncState;
output	[7:0]	HP2fp_L1RxUsr8B10BDispErr;
output	[11:0]	HP2fp_L1RxUsr8B10BEBCorCnt;
output	[11:0]	HP2fp_L1RxUsr8B10BEBStat;
output	[7:0]	HP2fp_L1RxUsr8B10BIsComma;
output	[7:0]	HP2fp_L1RxUsr8B10BIsK;
output	[7:0]	HP2fp_L1RxUsr8B10BNotInTable;
output	[7:0]	HP2fp_L1RxUsr8B10BRunDisp;
output	[0:0]	HP2fp_L1RxUsr8B10BValid;
output	[79:0]	HP2fp_L1RxUsrData;
output	[2:0]	HP2fp_L1RxUsrGBHeader;
output	[0:0]	HP2fp_L1RxUsrGBHeaderValid;
output	[0:0]	HP2fp_L1RxUsrGBStartSeq;
output	[2:0]	HP2fp_L1TxBufStatus;
output	[0:0]	HP2fp_L1TxSATAOOBComFinish;
output	[0:0]	HP2fp_L1TxUsrGBReady;
output	[0:0]	HP2fp_L0RxCALDetected;
output	[0:0]	HP2fp_L0RxGearboxIsSync;
output	[0:0]	HP2fp_L0RxOOBCOMINITDet;
output	[0:0]	HP2fp_L0RxOOBCOMSASDet;
output	[0:0]	HP2fp_L0RxOOBCOMWAKEDet;
output	[0:0]	HP2fp_L0RxOOBElecIdle;
output	[0:0]	HP2fp_L0RxOvrsmplErr;
output	[0:0]	HP2fp_L0RxPIPEPHYStatusRxDet;
output	[0:0]	HP2fp_L0RxPIPERxDetected;
output	[15:0]	HP2fp_L0RxPRBSErrCnt;
output	[15:0]	HP2fp_L0RxPRBSZeroCnt;
output	[1:0]	HP2fp_L0RxSyncState;
output	[7:0]	HP2fp_L0RxUsr8B10BDispErr;
output	[11:0]	HP2fp_L0RxUsr8B10BEBCorCnt;
output	[11:0]	HP2fp_L0RxUsr8B10BEBStat;
output	[7:0]	HP2fp_L0RxUsr8B10BIsComma;
output	[7:0]	HP2fp_L0RxUsr8B10BIsK;
output	[7:0]	HP2fp_L0RxUsr8B10BNotInTable;
output	[7:0]	HP2fp_L0RxUsr8B10BRunDisp;
output	[0:0]	HP2fp_L0RxUsr8B10BValid;
output	[79:0]	HP2fp_L0RxUsrData;
output	[2:0]	HP2fp_L0RxUsrGBHeader;
output	[0:0]	HP2fp_L0RxUsrGBHeaderValid;
output	[0:0]	HP2fp_L0RxUsrGBStartSeq;
output	[2:0]	HP2fp_L0TxBufStatus;
output	[0:0]	HP2fp_L0TxSATAOOBComFinish;
output	[0:0]	HP2fp_L0TxUsrGBReady;
output	[0:0]	HP2fp_PIPEPhyStatusForce;
output	[0:0]	HP2fp_PIPEPhyStatusSoft;
output	[0:0]	HP2fp_PowerOnDone;
output	[0:0]	HP2fp_RxLDuAlignAcqr;
output		HP2fp_xPLL_lockdet;
output		TSTCK3;
output		TSTCK2;
output		TSTCK1;
output		TSTCK0;
output		TXN3;
output		TXN2;
output		TXN1;
output		TXN0;
output		TXP3;
output		TXP2;
output		TXP1;
output		TXP0;
output		pbus_gnt;
output	[31:0]	pbus_rdata;
input		REFCLKN;
input		REFCLKP;
input		RXN3;
input		RXN2;
input		RXN1;
input		RXN0;
input		RXP3;
input		RXP2;
input		RXP1;
input		RXP0;
input		SP2HP_L3RXClkCorUse;
input		SP2HP_L3Rx8B10BDecMComDet;
input		SP2HP_L3Rx8B10BDecPComDet;
input		SP2HP_L3Rx8B10BUse;
input	[9:0]	SP2HP_L3Rx8B10BUserDefCom;
input		SP2HP_L3Rx8B10BValidComOnly;
input		SP2HP_L3Rx4B5BAlignEn;
input	[9:0]	SP2HP_L3Rx4B5BED;
input	[9:0]	SP2HP_L3Rx4B5BSD;
input		SP2HP_L3Rx4B5BUse;
input		SP2HP_L3RxBitReverse;
input		SP2HP_L3RxBufClr;
input	[1:0]	SP2HP_L3RxBufDepth;
input		SP2HP_L3RxBufUse;
input	[9:0]	SP2HP_L3RxCAL10BEnable;
input		SP2HP_L3RxCALAlignWord;
input		SP2HP_L3RxCALDetUse;
input		SP2HP_L3RxCALDouble;
input		SP2HP_L3RxCALEnMComAlign;
input		SP2HP_L3RxCALEnPComAlign;
input		SP2HP_L3RxCALMComDet;
input	[9:0]	SP2HP_L3RxCALMComValue;
input		SP2HP_L3RxCALPComDet;
input	[9:0]	SP2HP_L3RxCALPComValue;
input		SP2HP_L3RxCALSlide;
input	[1:0]	SP2HP_L3RxCALSlideMode;
input	[35:0]	SP2HP_L3RxCHBondSeq1;
input	[3:0]	SP2HP_L3RxCHBondSeq1En;
input	[8:0]	SP2HP_L3RxCHBondSeq1Mask;
input	[1:0]	SP2HP_L3RxClkCorAdjLen;
input	[8:0]	SP2HP_L3RxClkCorSeq14;
input	[8:0]	SP2HP_L3RxClkCorSeq13;
input	[8:0]	SP2HP_L3RxClkCorSeq12;
input	[8:0]	SP2HP_L3RxClkCorSeq11;
input	[3:0]	SP2HP_L3RxClkCorSeq1En;
input	[1:0]	SP2HP_L3RxDataWidth;
input		SP2HP_L3RxGearboxADJSel;
input		SP2HP_L3RxGearboxEnDec;
input		SP2HP_L3RxGearboxSlip;
input		SP2HP_L3RxGearboxUse;
input		SP2HP_L3RxInternalWidth;
input		SP2HP_L3RxLDEn;
input	[1:0]	SP2HP_L3RxNELClkMuxSel;
input	[1:0]	SP2HP_L3RxNLMux;
input		SP2HP_L3RxNLMuxWidth;
input	[2:0]	SP2HP_L3RxOOBBurstVal;
input	[5:0]	SP2HP_L3RxOOBMaxBurst;
input	[5:0]	SP2HP_L3RxOOBMaxCOMINIT;
input	[6:0]	SP2HP_L3RxOOBMaxCOMSAS;
input	[5:0]	SP2HP_L3RxOOBMaxCOMWAKE;
input	[5:0]	SP2HP_L3RxOOBMinBurst;
input	[5:0]	SP2HP_L3RxOOBMinCOMINIT;
input	[6:0]	SP2HP_L3RxOOBMinCOMSAS;
input	[5:0]	SP2HP_L3RxOOBMinCOMWAKE;
input		SP2HP_L3RxOvrsmplEnAlign;
input		SP2HP_L3RxOvrsmplMode;
input	[1:0]	SP2HP_L3RxPMux;
input		SP2HP_L3RxPRBSCntClr;
input	[2:0]	SP2HP_L3RxPRBSTst;
input	[39:0]	SP2HP_L3RxPRBSUsr;
input		SP2HP_L3RxPRBSWidth;
input		SP2HP_L3RxPRBSZCntClr;
input		SP2HP_L3RxPolarity;
input		SP2HP_L3RxRecClkMuxSel;
input		SP2HP_L3RxSyncEn;
input	[2:0]	SP2HP_L3RxSyncInvalidIncr;
input	[1:0]	SP2HP_L3RxSyncThres;
input	[2:0]	SP2HP_L3RxSyncThreshold;
input	[2:0]	SP2HP_L3RxUClk2MuxSel;
input	[1:0]	SP2HP_L3RxUClkMuxSel;
input		SP2HP_L3RxUsrClk;
input		SP2HP_L3RxUsrClk2;
input		SP2HP_L3Tx8B10BUse;
input		SP2HP_L3Tx4B5BUse;
input		SP2HP_L3TxBitReverse;
input		SP2HP_L3TxBufClr;
input		SP2HP_L3TxBufWidth;
input		SP2HP_L3TxBufferUse;
input	[1:0]	SP2HP_L3TxDMux;
input	[1:0]	SP2HP_L3TxDataWidth;
input		SP2HP_L3TxElecIdleAdj;
input	[1:0]	SP2HP_L3TxFlMux;
input	[1:0]	SP2HP_L3TxGearboxFunc;
input	[2:0]	SP2HP_L3TxGearboxReadyPre;
input		SP2HP_L3TxGearboxUse;
input		SP2HP_L3TxInternalWidth;
input	[1:0]	SP2HP_L3TxOOBMode;
input	[1:0]	SP2HP_L3TxOutClkMuxSel;
input		SP2HP_L3TxOvrsmplMode;
input	[1:0]	SP2HP_L3TxPCIEBeaconPWidth;
input		SP2HP_L3TxPCIEDetectRx;
input		SP2HP_L3TxPCIEElecIdle;
input		SP2HP_L3TxPClkMuxSel;
input	[2:0]	SP2HP_L3TxPMux;
input		SP2HP_L3TxPRBSErrCont;
input		SP2HP_L3TxPRBSErrOne;
input	[2:0]	SP2HP_L3TxPRBSTst;
input	[39:0]	SP2HP_L3TxPRBSUsr;
input		SP2HP_L3TxPRBSWidth;
input		SP2HP_L3TxPolarity;
input	[3:0]	SP2HP_L3TxSATAOOBComBurstVal;
input		SP2HP_L3TxSATAOOBComRESET;
input		SP2HP_L3TxSATAOOBComSAS;
input		SP2HP_L3TxSATAOOBComWAKE;
input		SP2HP_L3TxSATAOOBType;
input	[1:0]	SP2HP_L3TxUClk2MuxSel;
input	[1:0]	SP2HP_L3TxUClkMuxSel;
input	[1:0]	SP2HP_L3TxUIASmpl;
input	[7:0]	SP2HP_L3TxUsr8B10BDataK;
input	[7:0]	SP2HP_L3TxUsr8B10BDispMode;
input	[7:0]	SP2HP_L3TxUsr8B10BDispVal;
input		SP2HP_L3TxUsrClk;
input		SP2HP_L3TxUsrClk2;
input	[79:0]	SP2HP_L3TxUsrData;
input	[2:0]	SP2HP_L3TxUsrGBHeader;
input	[6:0]	SP2HP_L3TxUsrGBSequence;
input		SP2HP_L3TxUsrGBStartSeq;
input		SP2HP_L2RXClkCorUse;
input		SP2HP_L2Rx8B10BDecMComDet;
input		SP2HP_L2Rx8B10BDecPComDet;
input		SP2HP_L2Rx8B10BUse;
input	[9:0]	SP2HP_L2Rx8B10BUserDefCom;
input		SP2HP_L2Rx8B10BValidComOnly;
input		SP2HP_L2Rx4B5BAlignEn;
input	[9:0]	SP2HP_L2Rx4B5BED;
input	[9:0]	SP2HP_L2Rx4B5BSD;
input		SP2HP_L2Rx4B5BUse;
input		SP2HP_L2RxBitReverse;
input		SP2HP_L2RxBufClr;
input	[1:0]	SP2HP_L2RxBufDepth;
input		SP2HP_L2RxBufUse;
input	[9:0]	SP2HP_L2RxCAL10BEnable;
input		SP2HP_L2RxCALAlignWord;
input		SP2HP_L2RxCALDetUse;
input		SP2HP_L2RxCALDouble;
input		SP2HP_L2RxCALEnMComAlign;
input		SP2HP_L2RxCALEnPComAlign;
input		SP2HP_L2RxCALMComDet;
input	[9:0]	SP2HP_L2RxCALMComValue;
input		SP2HP_L2RxCALPComDet;
input	[9:0]	SP2HP_L2RxCALPComValue;
input		SP2HP_L2RxCALSlide;
input	[1:0]	SP2HP_L2RxCALSlideMode;
input	[35:0]	SP2HP_L2RxCHBondSeq1;
input	[3:0]	SP2HP_L2RxCHBondSeq1En;
input	[8:0]	SP2HP_L2RxCHBondSeq1Mask;
input	[1:0]	SP2HP_L2RxClkCorAdjLen;
input	[8:0]	SP2HP_L2RxClkCorSeq14;
input	[8:0]	SP2HP_L2RxClkCorSeq13;
input	[8:0]	SP2HP_L2RxClkCorSeq12;
input	[8:0]	SP2HP_L2RxClkCorSeq11;
input	[3:0]	SP2HP_L2RxClkCorSeq1En;
input	[1:0]	SP2HP_L2RxDataWidth;
input		SP2HP_L2RxGearboxADJSel;
input		SP2HP_L2RxGearboxEnDec;
input		SP2HP_L2RxGearboxSlip;
input		SP2HP_L2RxGearboxUse;
input		SP2HP_L2RxInternalWidth;
input		SP2HP_L2RxLDEn;
input	[1:0]	SP2HP_L2RxNELClkMuxSel;
input	[1:0]	SP2HP_L2RxNLMux;
input		SP2HP_L2RxNLMuxWidth;
input	[2:0]	SP2HP_L2RxOOBBurstVal;
input	[5:0]	SP2HP_L2RxOOBMaxBurst;
input	[5:0]	SP2HP_L2RxOOBMaxCOMINIT;
input	[6:0]	SP2HP_L2RxOOBMaxCOMSAS;
input	[5:0]	SP2HP_L2RxOOBMaxCOMWAKE;
input	[5:0]	SP2HP_L2RxOOBMinBurst;
input	[5:0]	SP2HP_L2RxOOBMinCOMINIT;
input	[6:0]	SP2HP_L2RxOOBMinCOMSAS;
input	[5:0]	SP2HP_L2RxOOBMinCOMWAKE;
input		SP2HP_L2RxOvrsmplEnAlign;
input		SP2HP_L2RxOvrsmplMode;
input	[1:0]	SP2HP_L2RxPMux;
input		SP2HP_L2RxPRBSCntClr;
input	[2:0]	SP2HP_L2RxPRBSTst;
input	[39:0]	SP2HP_L2RxPRBSUsr;
input		SP2HP_L2RxPRBSWidth;
input		SP2HP_L2RxPRBSZCntClr;
input		SP2HP_L2RxPolarity;
input		SP2HP_L2RxRecClkMuxSel;
input		SP2HP_L2RxSyncEn;
input	[2:0]	SP2HP_L2RxSyncInvalidIncr;
input	[1:0]	SP2HP_L2RxSyncThres;
input	[2:0]	SP2HP_L2RxSyncThreshold;
input	[2:0]	SP2HP_L2RxUClk2MuxSel;
input	[1:0]	SP2HP_L2RxUClkMuxSel;
input		SP2HP_L2RxUsrClk;
input		SP2HP_L2RxUsrClk2;
input		SP2HP_L2Tx8B10BUse;
input		SP2HP_L2Tx4B5BUse;
input		SP2HP_L2TxBitReverse;
input		SP2HP_L2TxBufClr;
input		SP2HP_L2TxBufWidth;
input		SP2HP_L2TxBufferUse;
input	[1:0]	SP2HP_L2TxDMux;
input	[1:0]	SP2HP_L2TxDataWidth;
input		SP2HP_L2TxElecIdleAdj;
input	[1:0]	SP2HP_L2TxFlMux;
input	[1:0]	SP2HP_L2TxGearboxFunc;
input	[2:0]	SP2HP_L2TxGearboxReadyPre;
input		SP2HP_L2TxGearboxUse;
input		SP2HP_L2TxInternalWidth;
input	[1:0]	SP2HP_L2TxOOBMode;
input	[1:0]	SP2HP_L2TxOutClkMuxSel;
input		SP2HP_L2TxOvrsmplMode;
input	[1:0]	SP2HP_L2TxPCIEBeaconPWidth;
input		SP2HP_L2TxPCIEDetectRx;
input		SP2HP_L2TxPCIEElecIdle;
input		SP2HP_L2TxPClkMuxSel;
input	[2:0]	SP2HP_L2TxPMux;
input		SP2HP_L2TxPRBSErrCont;
input		SP2HP_L2TxPRBSErrOne;
input	[2:0]	SP2HP_L2TxPRBSTst;
input	[39:0]	SP2HP_L2TxPRBSUsr;
input		SP2HP_L2TxPRBSWidth;
input		SP2HP_L2TxPolarity;
input	[3:0]	SP2HP_L2TxSATAOOBComBurstVal;
input		SP2HP_L2TxSATAOOBComRESET;
input		SP2HP_L2TxSATAOOBComSAS;
input		SP2HP_L2TxSATAOOBComWAKE;
input		SP2HP_L2TxSATAOOBType;
input	[1:0]	SP2HP_L2TxUClk2MuxSel;
input	[1:0]	SP2HP_L2TxUClkMuxSel;
input	[1:0]	SP2HP_L2TxUIASmpl;
input	[7:0]	SP2HP_L2TxUsr8B10BDataK;
input	[7:0]	SP2HP_L2TxUsr8B10BDispMode;
input	[7:0]	SP2HP_L2TxUsr8B10BDispVal;
input		SP2HP_L2TxUsrClk;
input		SP2HP_L2TxUsrClk2;
input	[79:0]	SP2HP_L2TxUsrData;
input	[2:0]	SP2HP_L2TxUsrGBHeader;
input	[6:0]	SP2HP_L2TxUsrGBSequence;
input		SP2HP_L2TxUsrGBStartSeq;
input		SP2HP_L1RXClkCorUse;
input		SP2HP_L1Rx8B10BDecMComDet;
input		SP2HP_L1Rx8B10BDecPComDet;
input		SP2HP_L1Rx8B10BUse;
input	[9:0]	SP2HP_L1Rx8B10BUserDefCom;
input		SP2HP_L1Rx8B10BValidComOnly;
input		SP2HP_L1Rx4B5BAlignEn;
input	[9:0]	SP2HP_L1Rx4B5BED;
input	[9:0]	SP2HP_L1Rx4B5BSD;
input		SP2HP_L1Rx4B5BUse;
input		SP2HP_L1RxBitReverse;
input		SP2HP_L1RxBufClr;
input	[1:0]	SP2HP_L1RxBufDepth;
input		SP2HP_L1RxBufUse;
input	[9:0]	SP2HP_L1RxCAL10BEnable;
input		SP2HP_L1RxCALAlignWord;
input		SP2HP_L1RxCALDetUse;
input		SP2HP_L1RxCALDouble;
input		SP2HP_L1RxCALEnMComAlign;
input		SP2HP_L1RxCALEnPComAlign;
input		SP2HP_L1RxCALMComDet;
input	[9:0]	SP2HP_L1RxCALMComValue;
input		SP2HP_L1RxCALPComDet;
input	[9:0]	SP2HP_L1RxCALPComValue;
input		SP2HP_L1RxCALSlide;
input	[1:0]	SP2HP_L1RxCALSlideMode;
input	[35:0]	SP2HP_L1RxCHBondSeq1;
input	[3:0]	SP2HP_L1RxCHBondSeq1En;
input	[8:0]	SP2HP_L1RxCHBondSeq1Mask;
input	[1:0]	SP2HP_L1RxClkCorAdjLen;
input	[8:0]	SP2HP_L1RxClkCorSeq14;
input	[8:0]	SP2HP_L1RxClkCorSeq13;
input	[8:0]	SP2HP_L1RxClkCorSeq12;
input	[8:0]	SP2HP_L1RxClkCorSeq11;
input	[3:0]	SP2HP_L1RxClkCorSeq1En;
input	[1:0]	SP2HP_L1RxDataWidth;
input		SP2HP_L1RxGearboxADJSel;
input		SP2HP_L1RxGearboxEnDec;
input		SP2HP_L1RxGearboxSlip;
input		SP2HP_L1RxGearboxUse;
input		SP2HP_L1RxInternalWidth;
input		SP2HP_L1RxLDEn;
input	[1:0]	SP2HP_L1RxNELClkMuxSel;
input	[1:0]	SP2HP_L1RxNLMux;
input		SP2HP_L1RxNLMuxWidth;
input	[2:0]	SP2HP_L1RxOOBBurstVal;
input	[5:0]	SP2HP_L1RxOOBMaxBurst;
input	[5:0]	SP2HP_L1RxOOBMaxCOMINIT;
input	[6:0]	SP2HP_L1RxOOBMaxCOMSAS;
input	[5:0]	SP2HP_L1RxOOBMaxCOMWAKE;
input	[5:0]	SP2HP_L1RxOOBMinBurst;
input	[5:0]	SP2HP_L1RxOOBMinCOMINIT;
input	[6:0]	SP2HP_L1RxOOBMinCOMSAS;
input	[5:0]	SP2HP_L1RxOOBMinCOMWAKE;
input		SP2HP_L1RxOvrsmplEnAlign;
input		SP2HP_L1RxOvrsmplMode;
input	[1:0]	SP2HP_L1RxPMux;
input		SP2HP_L1RxPRBSCntClr;
input	[2:0]	SP2HP_L1RxPRBSTst;
input	[39:0]	SP2HP_L1RxPRBSUsr;
input		SP2HP_L1RxPRBSWidth;
input		SP2HP_L1RxPRBSZCntClr;
input		SP2HP_L1RxPolarity;
input		SP2HP_L1RxRecClkMuxSel;
input		SP2HP_L1RxSyncEn;
input	[2:0]	SP2HP_L1RxSyncInvalidIncr;
input	[1:0]	SP2HP_L1RxSyncThres;
input	[2:0]	SP2HP_L1RxSyncThreshold;
input	[2:0]	SP2HP_L1RxUClk2MuxSel;
input	[1:0]	SP2HP_L1RxUClkMuxSel;
input		SP2HP_L1RxUsrClk;
input		SP2HP_L1RxUsrClk2;
input		SP2HP_L1Tx8B10BUse;
input		SP2HP_L1Tx4B5BUse;
input		SP2HP_L1TxBitReverse;
input		SP2HP_L1TxBufClr;
input		SP2HP_L1TxBufWidth;
input		SP2HP_L1TxBufferUse;
input	[1:0]	SP2HP_L1TxDMux;
input	[1:0]	SP2HP_L1TxDataWidth;
input		SP2HP_L1TxElecIdleAdj;
input	[1:0]	SP2HP_L1TxFlMux;
input	[1:0]	SP2HP_L1TxGearboxFunc;
input	[2:0]	SP2HP_L1TxGearboxReadyPre;
input		SP2HP_L1TxGearboxUse;
input		SP2HP_L1TxInternalWidth;
input	[1:0]	SP2HP_L1TxOOBMode;
input	[1:0]	SP2HP_L1TxOutClkMuxSel;
input		SP2HP_L1TxOvrsmplMode;
input	[1:0]	SP2HP_L1TxPCIEBeaconPWidth;
input		SP2HP_L1TxPCIEDetectRx;
input		SP2HP_L1TxPCIEElecIdle;
input		SP2HP_L1TxPClkMuxSel;
input	[2:0]	SP2HP_L1TxPMux;
input		SP2HP_L1TxPRBSErrCont;
input		SP2HP_L1TxPRBSErrOne;
input	[2:0]	SP2HP_L1TxPRBSTst;
input	[39:0]	SP2HP_L1TxPRBSUsr;
input		SP2HP_L1TxPRBSWidth;
input		SP2HP_L1TxPolarity;
input	[3:0]	SP2HP_L1TxSATAOOBComBurstVal;
input		SP2HP_L1TxSATAOOBComRESET;
input		SP2HP_L1TxSATAOOBComSAS;
input		SP2HP_L1TxSATAOOBComWAKE;
input		SP2HP_L1TxSATAOOBType;
input	[1:0]	SP2HP_L1TxUClk2MuxSel;
input	[1:0]	SP2HP_L1TxUClkMuxSel;
input	[1:0]	SP2HP_L1TxUIASmpl;
input	[7:0]	SP2HP_L1TxUsr8B10BDataK;
input	[7:0]	SP2HP_L1TxUsr8B10BDispMode;
input	[7:0]	SP2HP_L1TxUsr8B10BDispVal;
input		SP2HP_L1TxUsrClk;
input		SP2HP_L1TxUsrClk2;
input	[79:0]	SP2HP_L1TxUsrData;
input	[2:0]	SP2HP_L1TxUsrGBHeader;
input	[6:0]	SP2HP_L1TxUsrGBSequence;
input		SP2HP_L1TxUsrGBStartSeq;
input		SP2HP_L0RXClkCorUse;
input		SP2HP_L0Rx8B10BDecMComDet;
input		SP2HP_L0Rx8B10BDecPComDet;
input		SP2HP_L0Rx8B10BUse;
input	[9:0]	SP2HP_L0Rx8B10BUserDefCom;
input		SP2HP_L0Rx8B10BValidComOnly;
input		SP2HP_L0Rx4B5BAlignEn;
input	[9:0]	SP2HP_L0Rx4B5BED;
input	[9:0]	SP2HP_L0Rx4B5BSD;
input		SP2HP_L0Rx4B5BUse;
input		SP2HP_L0RxBitReverse;
input		SP2HP_L0RxBufClr;
input	[1:0]	SP2HP_L0RxBufDepth;
input		SP2HP_L0RxBufUse;
input	[9:0]	SP2HP_L0RxCAL10BEnable;
input		SP2HP_L0RxCALAlignWord;
input		SP2HP_L0RxCALDetUse;
input		SP2HP_L0RxCALDouble;
input		SP2HP_L0RxCALEnMComAlign;
input		SP2HP_L0RxCALEnPComAlign;
input		SP2HP_L0RxCALMComDet;
input	[9:0]	SP2HP_L0RxCALMComValue;
input		SP2HP_L0RxCALPComDet;
input	[9:0]	SP2HP_L0RxCALPComValue;
input		SP2HP_L0RxCALSlide;
input	[1:0]	SP2HP_L0RxCALSlideMode;
input	[35:0]	SP2HP_L0RxCHBondSeq1;
input	[3:0]	SP2HP_L0RxCHBondSeq1En;
input	[8:0]	SP2HP_L0RxCHBondSeq1Mask;
input	[1:0]	SP2HP_L0RxClkCorAdjLen;
input	[8:0]	SP2HP_L0RxClkCorSeq14;
input	[8:0]	SP2HP_L0RxClkCorSeq13;
input	[8:0]	SP2HP_L0RxClkCorSeq12;
input	[8:0]	SP2HP_L0RxClkCorSeq11;
input	[3:0]	SP2HP_L0RxClkCorSeq1En;
input	[1:0]	SP2HP_L0RxDataWidth;
input		SP2HP_L0RxGearboxADJSel;
input		SP2HP_L0RxGearboxEnDec;
input		SP2HP_L0RxGearboxSlip;
input		SP2HP_L0RxGearboxUse;
input		SP2HP_L0RxInternalWidth;
input		SP2HP_L0RxLDEn;
input	[1:0]	SP2HP_L0RxNELClkMuxSel;
input	[1:0]	SP2HP_L0RxNLMux;
input		SP2HP_L0RxNLMuxWidth;
input	[2:0]	SP2HP_L0RxOOBBurstVal;
input	[5:0]	SP2HP_L0RxOOBMaxBurst;
input	[5:0]	SP2HP_L0RxOOBMaxCOMINIT;
input	[6:0]	SP2HP_L0RxOOBMaxCOMSAS;
input	[5:0]	SP2HP_L0RxOOBMaxCOMWAKE;
input	[5:0]	SP2HP_L0RxOOBMinBurst;
input	[5:0]	SP2HP_L0RxOOBMinCOMINIT;
input	[6:0]	SP2HP_L0RxOOBMinCOMSAS;
input	[5:0]	SP2HP_L0RxOOBMinCOMWAKE;
input		SP2HP_L0RxOvrsmplEnAlign;
input		SP2HP_L0RxOvrsmplMode;
input	[1:0]	SP2HP_L0RxPMux;
input		SP2HP_L0RxPRBSCntClr;
input	[2:0]	SP2HP_L0RxPRBSTst;
input	[39:0]	SP2HP_L0RxPRBSUsr;
input		SP2HP_L0RxPRBSWidth;
input		SP2HP_L0RxPRBSZCntClr;
input		SP2HP_L0RxPolarity;
input		SP2HP_L0RxRecClkMuxSel;
input		SP2HP_L0RxSyncEn;
input	[2:0]	SP2HP_L0RxSyncInvalidIncr;
input	[1:0]	SP2HP_L0RxSyncThres;
input	[2:0]	SP2HP_L0RxSyncThreshold;
input	[2:0]	SP2HP_L0RxUClk2MuxSel;
input	[1:0]	SP2HP_L0RxUClkMuxSel;
input		SP2HP_L0RxUsrClk;
input		SP2HP_L0RxUsrClk2;
input		SP2HP_L0Tx8B10BUse;
input		SP2HP_L0Tx4B5BUse;
input		SP2HP_L0TxBitReverse;
input		SP2HP_L0TxBufClr;
input		SP2HP_L0TxBufWidth;
input		SP2HP_L0TxBufferUse;
input	[1:0]	SP2HP_L0TxDMux;
input	[1:0]	SP2HP_L0TxDataWidth;
input		SP2HP_L0TxElecIdleAdj;
input	[1:0]	SP2HP_L0TxFlMux;
input	[1:0]	SP2HP_L0TxGearboxFunc;
input	[2:0]	SP2HP_L0TxGearboxReadyPre;
input		SP2HP_L0TxGearboxUse;
input		SP2HP_L0TxInternalWidth;
input	[1:0]	SP2HP_L0TxOOBMode;
input	[1:0]	SP2HP_L0TxOutClkMuxSel;
input		SP2HP_L0TxOvrsmplMode;
input	[1:0]	SP2HP_L0TxPCIEBeaconPWidth;
input		SP2HP_L0TxPCIEDetectRx;
input		SP2HP_L0TxPCIEElecIdle;
input		SP2HP_L0TxPClkMuxSel;
input	[2:0]	SP2HP_L0TxPMux;
input		SP2HP_L0TxPRBSErrCont;
input		SP2HP_L0TxPRBSErrOne;
input	[2:0]	SP2HP_L0TxPRBSTst;
input	[39:0]	SP2HP_L0TxPRBSUsr;
input		SP2HP_L0TxPRBSWidth;
input		SP2HP_L0TxPolarity;
input	[3:0]	SP2HP_L0TxSATAOOBComBurstVal;
input		SP2HP_L0TxSATAOOBComRESET;
input		SP2HP_L0TxSATAOOBComSAS;
input		SP2HP_L0TxSATAOOBComWAKE;
input		SP2HP_L0TxSATAOOBType;
input	[1:0]	SP2HP_L0TxUClk2MuxSel;
input	[1:0]	SP2HP_L0TxUClkMuxSel;
input	[1:0]	SP2HP_L0TxUIASmpl;
input	[7:0]	SP2HP_L0TxUsr8B10BDataK;
input	[7:0]	SP2HP_L0TxUsr8B10BDispMode;
input	[7:0]	SP2HP_L0TxUsr8B10BDispVal;
input		SP2HP_L0TxUsrClk;
input		SP2HP_L0TxUsrClk2;
input	[79:0]	SP2HP_L0TxUsrData;
input	[2:0]	SP2HP_L0TxUsrGBHeader;
input	[6:0]	SP2HP_L0TxUsrGBSequence;
input		SP2HP_L0TxUsrGBStartSeq;
input	[3:0]	SP2HP_LaneEn;
input	[1:0]	SP2HP_PCIEMode;
input	[13:0]	SP2HP_PonChgClkT2;
input	[13:0]	SP2HP_PonChgClkT1;
input	[13:0]	SP2HP_PonDfeCalT;
input	[13:0]	SP2HP_PonInitT;
input	[13:0]	SP2HP_PonOfstCalHiT;
input	[13:0]	SP2HP_PonOfstCalLoT;
input	[13:0]	SP2HP_PonPllDetT;
input	[13:0]	SP2HP_PonPreDfeCalT;
input	[13:0]	SP2HP_PonPrePllDetT;
input	[13:0]	SP2HP_PonPreResCalT;
input	[13:0]	SP2HP_PonPwrIntvalT;
input	[13:0]	SP2HP_PonResCalHiT;
input	[13:0]	SP2HP_PonResCalLoT;
input	[3:0]	SP2HP_RxUnifClkSel;
input		SP2HP_RxX4Mode;
input		SP2HP_SSCEnX4;
input		SP2HP_SysRstBSel;
input	[6:0]	SP2HP_TxDetRxT4;
input	[2:0]	SP2HP_TxDetRxT3;
input	[2:0]	SP2HP_TxDetRxT2;
input	[5:0]	SP2HP_TxDetRxT1;
input	[13:0]	SP2HP_TxPhaseAlignT;
input		SP2HP_TxX4Mode;
input		SP2HP_UsrRst_N;
input		SP2HP_UsrRxRst_N;
input		SP2HP_UsrTxRst_N;
input		SP2HP_xBG_SafeMode;
input	[3:0]	SP2HP_xBG_pr200clkmux;
input	[3:0]	SP2HP_xBG_pr100BRCal;
input	[3:0]	SP2HP_xBG_pr100Rx;
input	[3:0]	SP2HP_xBG_pr100Tx;
input	[3:0]	SP2HP_xBG_pr100spare;
input	[3:0]	SP2HP_xBG_prcal100Rx;
input	[3:0]	SP2HP_xBG_prcal100Tx;
input	[1:0]	SP2HP_xBG_prcal50Pll;
input	[1:0]	SP2HP_xBG_prcal50spare;
input		SP2HP_xBG_pwrdnB;
input	[2:0]	SP2HP_xBG_trim;
input	[1:0]	SP2HP_xCDR3_PIbiasTrim;
input	[2:0]	SP2HP_xCDR3_PIcapTrim;
input	[1:0]	SP2HP_xCDR3_PdivSelRx;
input		SP2HP_xCDR3_SelFourFive;
input		SP2HP_xCDR3_clkmode;
input		SP2HP_xCDR3_dccen;
input		SP2HP_xCDR3_dccfix;
input		SP2HP_xCDR3_dcctrim;
input		SP2HP_xCDR3_hold;
input	[3:0]	SP2HP_xCDR3_inc;
input	[4:0]	SP2HP_xCDR3_incF;
input	[4:0]	SP2HP_xCDR3_limHF;
input	[4:0]	SP2HP_xCDR3_limLF;
input		SP2HP_xCDR3_metamode;
input		SP2HP_xCDR3_mult2F;
input	[7:0]	SP2HP_xCDR3_offs;
input		SP2HP_xCDR3_pwrdnB;
input		SP2HP_xCDR3_updnsw;
input	[1:0]	SP2HP_xCDR2_PIbiasTrim;
input	[2:0]	SP2HP_xCDR2_PIcapTrim;
input	[1:0]	SP2HP_xCDR2_PdivSelRx;
input		SP2HP_xCDR2_SelFourFive;
input		SP2HP_xCDR2_clkmode;
input		SP2HP_xCDR2_dccen;
input		SP2HP_xCDR2_dccfix;
input		SP2HP_xCDR2_dcctrim;
input		SP2HP_xCDR2_hold;
input	[3:0]	SP2HP_xCDR2_inc;
input	[4:0]	SP2HP_xCDR2_incF;
input	[4:0]	SP2HP_xCDR2_limHF;
input	[4:0]	SP2HP_xCDR2_limLF;
input		SP2HP_xCDR2_metamode;
input		SP2HP_xCDR2_mult2F;
input	[7:0]	SP2HP_xCDR2_offs;
input		SP2HP_xCDR2_pwrdnB;
input		SP2HP_xCDR2_updnsw;
input	[1:0]	SP2HP_xCDR1_PIbiasTrim;
input	[2:0]	SP2HP_xCDR1_PIcapTrim;
input	[1:0]	SP2HP_xCDR1_PdivSelRx;
input		SP2HP_xCDR1_SelFourFive;
input		SP2HP_xCDR1_clkmode;
input		SP2HP_xCDR1_dccen;
input		SP2HP_xCDR1_dccfix;
input		SP2HP_xCDR1_dcctrim;
input		SP2HP_xCDR1_hold;
input	[3:0]	SP2HP_xCDR1_inc;
input	[4:0]	SP2HP_xCDR1_incF;
input	[4:0]	SP2HP_xCDR1_limHF;
input	[4:0]	SP2HP_xCDR1_limLF;
input		SP2HP_xCDR1_metamode;
input		SP2HP_xCDR1_mult2F;
input	[7:0]	SP2HP_xCDR1_offs;
input		SP2HP_xCDR1_pwrdnB;
input		SP2HP_xCDR1_updnsw;
input	[1:0]	SP2HP_xCDR0_PIbiasTrim;
input	[2:0]	SP2HP_xCDR0_PIcapTrim;
input	[1:0]	SP2HP_xCDR0_PdivSelRx;
input		SP2HP_xCDR0_SelFourFive;
input		SP2HP_xCDR0_clkmode;
input		SP2HP_xCDR0_dccen;
input		SP2HP_xCDR0_dccfix;
input		SP2HP_xCDR0_dcctrim;
input		SP2HP_xCDR0_hold;
input	[3:0]	SP2HP_xCDR0_inc;
input	[4:0]	SP2HP_xCDR0_incF;
input	[4:0]	SP2HP_xCDR0_limHF;
input	[4:0]	SP2HP_xCDR0_limLF;
input		SP2HP_xCDR0_metamode;
input		SP2HP_xCDR0_mult2F;
input	[7:0]	SP2HP_xCDR0_offs;
input		SP2HP_xCDR0_pwrdnB;
input		SP2HP_xCDR0_updnsw;
input		SP2HP_xCMU_clkmux_pwrdnB;
input		SP2HP_xCMU_clkmux_swon;
input	[1:0]	SP2HP_xCMU_cur_trim;
input		SP2HP_xCMU_pwrdnB;
input	[5:0]	SP2HP_xCMU_refclk_sel;
input		SP2HP_xCTLE3_Adaps_En;
input	[1:0]	SP2HP_xCTLE3_Adaps_inc;
input	[3:0]	SP2HP_xCTLE3_memCap;
input	[2:0]	SP2HP_xCTLE3_memRes3;
input	[1:0]	SP2HP_xCTLE3_memRes2;
input	[1:0]	SP2HP_xCTLE3_memRes1;
input		SP2HP_xCTLE2_Adaps_En;
input	[1:0]	SP2HP_xCTLE2_Adaps_inc;
input	[3:0]	SP2HP_xCTLE2_memCap;
input	[2:0]	SP2HP_xCTLE2_memRes3;
input	[1:0]	SP2HP_xCTLE2_memRes2;
input	[1:0]	SP2HP_xCTLE2_memRes1;
input		SP2HP_xCTLE1_Adaps_En;
input	[1:0]	SP2HP_xCTLE1_Adaps_inc;
input	[3:0]	SP2HP_xCTLE1_memCap;
input	[2:0]	SP2HP_xCTLE1_memRes3;
input	[1:0]	SP2HP_xCTLE1_memRes2;
input	[1:0]	SP2HP_xCTLE1_memRes1;
input		SP2HP_xCTLE0_Adaps_En;
input	[1:0]	SP2HP_xCTLE0_Adaps_inc;
input	[3:0]	SP2HP_xCTLE0_memCap;
input	[2:0]	SP2HP_xCTLE0_memRes3;
input	[1:0]	SP2HP_xCTLE0_memRes2;
input	[1:0]	SP2HP_xCTLE0_memRes1;
input		SP2HP_xDFE3_Adaps_En;
input		SP2HP_xDFE3_AnaClkEn;
input		SP2HP_xDFE3_EyeScan_En;
input	[4:0]	SP2HP_xDFE3_eqGain;
input	[2:0]	SP2HP_xDFE3_isoGain;
input	[5:0]	SP2HP_xDFE3_memDly;
input	[3:0]	SP2HP_xDFE3_memTap4;
input	[3:0]	SP2HP_xDFE3_memTap3;
input	[4:0]	SP2HP_xDFE3_memTap2;
input	[4:0]	SP2HP_xDFE3_memTap1;
input		SP2HP_xDFE3_setDly;
input		SP2HP_xDFE3_setEq;
input		SP2HP_xDFE3_tapcursel;
input		SP2HP_xDFE2_Adaps_En;
input		SP2HP_xDFE2_AnaClkEn;
input		SP2HP_xDFE2_EyeScan_En;
input	[4:0]	SP2HP_xDFE2_eqGain;
input	[2:0]	SP2HP_xDFE2_isoGain;
input	[5:0]	SP2HP_xDFE2_memDly;
input	[3:0]	SP2HP_xDFE2_memTap4;
input	[3:0]	SP2HP_xDFE2_memTap3;
input	[4:0]	SP2HP_xDFE2_memTap2;
input	[4:0]	SP2HP_xDFE2_memTap1;
input		SP2HP_xDFE2_setDly;
input		SP2HP_xDFE2_setEq;
input		SP2HP_xDFE2_tapcursel;
input		SP2HP_xDFE1_Adaps_En;
input		SP2HP_xDFE1_AnaClkEn;
input		SP2HP_xDFE1_EyeScan_En;
input	[4:0]	SP2HP_xDFE1_eqGain;
input	[2:0]	SP2HP_xDFE1_isoGain;
input	[5:0]	SP2HP_xDFE1_memDly;
input	[3:0]	SP2HP_xDFE1_memTap4;
input	[3:0]	SP2HP_xDFE1_memTap3;
input	[4:0]	SP2HP_xDFE1_memTap2;
input	[4:0]	SP2HP_xDFE1_memTap1;
input		SP2HP_xDFE1_setDly;
input		SP2HP_xDFE1_setEq;
input		SP2HP_xDFE1_tapcursel;
input		SP2HP_xDFE0_Adaps_En;
input		SP2HP_xDFE0_AnaClkEn;
input		SP2HP_xDFE0_EyeScan_En;
input	[4:0]	SP2HP_xDFE0_eqGain;
input	[2:0]	SP2HP_xDFE0_isoGain;
input	[5:0]	SP2HP_xDFE0_memDly;
input	[3:0]	SP2HP_xDFE0_memTap4;
input	[3:0]	SP2HP_xDFE0_memTap3;
input	[4:0]	SP2HP_xDFE0_memTap2;
input	[4:0]	SP2HP_xDFE0_memTap1;
input		SP2HP_xDFE0_setDly;
input		SP2HP_xDFE0_setEq;
input		SP2HP_xDFE0_tapcursel;
input		SP2HP_xDFECalEn3_mem;
input		SP2HP_xDFECalEn3_sel;
input		SP2HP_xDFECalEn2_mem;
input		SP2HP_xDFECalEn2_sel;
input		SP2HP_xDFECalEn1_mem;
input		SP2HP_xDFECalEn1_sel;
input		SP2HP_xDFECalEn0_mem;
input		SP2HP_xDFECalEn0_sel;
input		SP2HP_xJTAG_AC_Signal;
input		SP2HP_xJTAG_ClockDR;
input		SP2HP_xJTAG_En;
input		SP2HP_xJTAG_ShiftDR;
input		SP2HP_xJTAG_UpdateDR;
input		SP2HP_xJTAG_acmode;
input		SP2HP_xJTAG_ini_mem;
input		SP2HP_xJTAG_pwrdnB;
input		SP2HP_xJTAG_tap_resetB;
input		SP2HP_xJTAG_tdi;
input		SP2HP_xLane3_farlpbken;
input		SP2HP_xLane3_nearlpbken;
input		SP2HP_xLane2_farlpbken;
input		SP2HP_xLane2_nearlpbken;
input		SP2HP_xLane1_farlpbken;
input		SP2HP_xLane1_nearlpbken;
input		SP2HP_xLane0_farlpbken;
input		SP2HP_xLane0_nearlpbken;
input		SP2HP_xMisc_pwrdnB;
input		SP2HP_xMisc_resetB;
input		SP2HP_xOSC_CrntEn;
input		SP2HP_xOSC_FSEn;
input	[3:0]	SP2HP_xOSC_Rtrim;
input		SP2HP_xOSC_pwrdnB;
input		SP2HP_xOfstCal3_Ovrd;
input	[1:0]	SP2HP_xOfstCal3_inc;
input	[4:0]	SP2HP_xOfstCal3_mem;
input		SP2HP_xOfstCal3_memCtrl;
input		SP2HP_xOfstCal3_memEn;
input		SP2HP_xOfstCal3_pwrdnB;
input		SP2HP_xOfstCal2_Ovrd;
input	[1:0]	SP2HP_xOfstCal2_inc;
input	[4:0]	SP2HP_xOfstCal2_mem;
input		SP2HP_xOfstCal2_memCtrl;
input		SP2HP_xOfstCal2_memEn;
input		SP2HP_xOfstCal2_pwrdnB;
input		SP2HP_xOfstCal1_Ovrd;
input	[1:0]	SP2HP_xOfstCal1_inc;
input	[4:0]	SP2HP_xOfstCal1_mem;
input		SP2HP_xOfstCal1_memCtrl;
input		SP2HP_xOfstCal1_memEn;
input		SP2HP_xOfstCal1_pwrdnB;
input		SP2HP_xOfstCal0_Ovrd;
input	[1:0]	SP2HP_xOfstCal0_inc;
input	[4:0]	SP2HP_xOfstCal0_mem;
input		SP2HP_xOfstCal0_memCtrl;
input		SP2HP_xOfstCal0_memEn;
input		SP2HP_xOfstCal0_pwrdnB;
input		SP2HP_xPLL_CntlLimit_en;
input	[5:0]	SP2HP_xPLL_FBDIV;
input		SP2HP_xPLL_LockDet_Force_Lock;
input	[3:0]	SP2HP_xPLL_Qpump_2;
input	[3:0]	SP2HP_xPLL_Qpump_1;
input	[5:0]	SP2HP_xPLL_REFDIV;
input	[2:0]	SP2HP_xPLL_VCO_Ctuning;
input	[2:0]	SP2HP_xPLL_buf_Itrim;
input		SP2HP_xPLL_lockdet_en;
input	[1:0]	SP2HP_xPLL_lockdet_period_sel;
input	[2:0]	SP2HP_xPLL_lockdet_ppm_sel1;
input	[2:0]	SP2HP_xPLL_lockdet_ppm_sel0;
input	[1:0]	SP2HP_xPLL_pdivSel;
input		SP2HP_xPLL_pwrdnB;
input		SP2HP_xPLL_resetB;
input		SP2HP_xPLL_selFourFive;
input		SP2HP_xRX3_busdivSel;
input		SP2HP_xRX3_pwrdnB;
input		SP2HP_xRX3_set_phase;
input		SP2HP_xRX3_slip_clk;
input		SP2HP_xRX3_syncRxToUsrclk;
input		SP2HP_xRX3_xrChicoOvrPh5to9;
input	[4:0]	SP2HP_xRX3_xrChicoOvrd;
input		SP2HP_xRX3_xrChicoOvrdEn;
input		SP2HP_xRX2_busdivSel;
input		SP2HP_xRX2_pwrdnB;
input		SP2HP_xRX2_set_phase;
input		SP2HP_xRX2_slip_clk;
input		SP2HP_xRX2_syncRxToUsrclk;
input		SP2HP_xRX2_xrChicoOvrPh5to9;
input	[4:0]	SP2HP_xRX2_xrChicoOvrd;
input		SP2HP_xRX2_xrChicoOvrdEn;
input		SP2HP_xRX1_busdivSel;
input		SP2HP_xRX1_pwrdnB;
input		SP2HP_xRX1_set_phase;
input		SP2HP_xRX1_slip_clk;
input		SP2HP_xRX1_syncRxToUsrclk;
input		SP2HP_xRX1_xrChicoOvrPh5to9;
input	[4:0]	SP2HP_xRX1_xrChicoOvrd;
input		SP2HP_xRX1_xrChicoOvrdEn;
input		SP2HP_xRX0_busdivSel;
input		SP2HP_xRX0_pwrdnB;
input		SP2HP_xRX0_set_phase;
input		SP2HP_xRX0_slip_clk;
input		SP2HP_xRX0_syncRxToUsrclk;
input		SP2HP_xRX0_xrChicoOvrPh5to9;
input	[4:0]	SP2HP_xRX0_xrChicoOvrd;
input		SP2HP_xRX0_xrChicoOvrdEn;
input	[1:0]	SP2HP_xRXAFE3_InCMTrim;
input		SP2HP_xRXAFE3_rcvShuntEn;
input		SP2HP_xRXAFE3_rcvVssTermEn;
input		SP2HP_xRXAFE3_rcvVttTermEn;
input		SP2HP_xRXAFE3_termRes50En;
input	[1:0]	SP2HP_xRXAFE2_InCMTrim;
input		SP2HP_xRXAFE2_rcvShuntEn;
input		SP2HP_xRXAFE2_rcvVssTermEn;
input		SP2HP_xRXAFE2_rcvVttTermEn;
input		SP2HP_xRXAFE2_termRes50En;
input	[1:0]	SP2HP_xRXAFE1_InCMTrim;
input		SP2HP_xRXAFE1_rcvShuntEn;
input		SP2HP_xRXAFE1_rcvVssTermEn;
input		SP2HP_xRXAFE1_rcvVttTermEn;
input		SP2HP_xRXAFE1_termRes50En;
input	[1:0]	SP2HP_xRXAFE0_InCMTrim;
input		SP2HP_xRXAFE0_rcvShuntEn;
input		SP2HP_xRXAFE0_rcvVssTermEn;
input		SP2HP_xRXAFE0_rcvVttTermEn;
input		SP2HP_xRXAFE0_termRes50En;
input	[2:0]	SP2HP_xRXSquelch3_noSigLevel;
input		SP2HP_xRXSquelch3_pwrdnB;
input	[2:0]	SP2HP_xRXSquelch2_noSigLevel;
input		SP2HP_xRXSquelch2_pwrdnB;
input	[2:0]	SP2HP_xRXSquelch1_noSigLevel;
input		SP2HP_xRXSquelch1_pwrdnB;
input	[2:0]	SP2HP_xRXSquelch0_noSigLevel;
input		SP2HP_xRXSquelch0_pwrdnB;
input	[2:0]	SP2HP_xResCal_Bg_offset;
input	[2:0]	SP2HP_xResCal_LPF_offset;
input		SP2HP_xResCal_MemCtrl;
input		SP2HP_xResCal_MemEn;
input	[4:0]	SP2HP_xResCal_MemRes_Bg;
input	[4:0]	SP2HP_xResCal_MemRes_LPF;
input	[4:0]	SP2HP_xResCal_MemRes_Rx;
input	[4:0]	SP2HP_xResCal_MemRes_Tx;
input		SP2HP_xResCal_ResBg_sel;
input		SP2HP_xResCal_ResLPF_sel;
input		SP2HP_xResCal_ResRx_sel;
input		SP2HP_xResCal_ResTx_sel;
input	[2:0]	SP2HP_xResCal_Rx_offset;
input	[2:0]	SP2HP_xResCal_Tx_offset;
input	[4:0]	SP2HP_xTOP_DivOOB;
input	[4:0]	SP2HP_xTOP_DivSSC;
input	[4:0]	SP2HP_xTOP_DivSYS;
input		SP2HP_xTOP_SYSClkSel;
input		SP2HP_xTX3_ACCCLK_ROTATEH;
input		SP2HP_xTX3_ACC_DIN_SEL;
input	[1:0]	SP2HP_xTX3_ACC_NSEL;
input	[7:0]	SP2HP_xTX3_ACC_OVERRIDE;
input		SP2HP_xTX3_ACC_OVERRIDE_EN;
input		SP2HP_xTX3_ACC_ROTATE;
input		SP2HP_xTX3_ACC_UPDNSW;
input		SP2HP_xTX3_Clk_pwrdnB;
input	[2:0]	SP2HP_xTX3_DrvPostCursor;
input	[2:0]	SP2HP_xTX3_DrvPreCursor;
input		SP2HP_xTX3_Drv_pwrdnB;
input	[2:0]	SP2HP_xTX3_Drvbiastrim;
input	[3:0]	SP2HP_xTX3_Drvswing;
input	[2:0]	SP2HP_xTX3_PI_captrim;
input		SP2HP_xTX3_PI_pwrdnB;
input	[1:0]	SP2HP_xTX3_PIbiasTrim;
input		SP2HP_xTX3_Resl_En;
input		SP2HP_xTX3_SSC_EN;
input	[8:0]	SP2HP_xTX3_SSC_OVERRIDE;
input		SP2HP_xTX3_SSC_OVERRIDE_EN;
input	[4:0]	SP2HP_xTX3_SSC_TSEL;
input		SP2HP_xTX3_Ser_pwrdnB;
input	[2:0]	SP2HP_xTX3_Serbiastrim;
input	[3:0]	SP2HP_xTX3_Vreftrim;
input		SP2HP_xTX3_activepkEn;
input		SP2HP_xTX3_busdivSel;
input		SP2HP_xTX3_chico_cksel;
input		SP2HP_xTX3_chico_pwrdnB;
input	[2:0]	SP2HP_xTX3_ctune;
input	[1:0]	SP2HP_xTX3_dccbiastrim;
input	[1:0]	SP2HP_xTX3_dccerrtrim;
input		SP2HP_xTX3_dccfix;
input	[2:0]	SP2HP_xTX3_gmtune;
input		SP2HP_xTX3_ovsdivEn;
input	[1:0]	SP2HP_xTX3_pdivSel;
input		SP2HP_xTX3_pwrdnB;
input		SP2HP_xTX3_selFourFive;
input		SP2HP_xTX3_sendidle;
input		SP2HP_xTX3_syncTxToUsrclk;
input		SP2HP_xTX3_tdccEn;
input		SP2HP_xTX3_tdccovrd;
input		SP2HP_xTX2_ACCCLK_ROTATEH;
input		SP2HP_xTX2_ACC_DIN_SEL;
input	[1:0]	SP2HP_xTX2_ACC_NSEL;
input	[7:0]	SP2HP_xTX2_ACC_OVERRIDE;
input		SP2HP_xTX2_ACC_OVERRIDE_EN;
input		SP2HP_xTX2_ACC_ROTATE;
input		SP2HP_xTX2_ACC_UPDNSW;
input		SP2HP_xTX2_Clk_pwrdnB;
input	[2:0]	SP2HP_xTX2_DrvPostCursor;
input	[2:0]	SP2HP_xTX2_DrvPreCursor;
input		SP2HP_xTX2_Drv_pwrdnB;
input	[2:0]	SP2HP_xTX2_Drvbiastrim;
input	[3:0]	SP2HP_xTX2_Drvswing;
input	[2:0]	SP2HP_xTX2_PI_captrim;
input		SP2HP_xTX2_PI_pwrdnB;
input	[1:0]	SP2HP_xTX2_PIbiasTrim;
input		SP2HP_xTX2_Resl_En;
input		SP2HP_xTX2_SSC_EN;
input	[8:0]	SP2HP_xTX2_SSC_OVERRIDE;
input		SP2HP_xTX2_SSC_OVERRIDE_EN;
input	[4:0]	SP2HP_xTX2_SSC_TSEL;
input		SP2HP_xTX2_Ser_pwrdnB;
input	[2:0]	SP2HP_xTX2_Serbiastrim;
input	[3:0]	SP2HP_xTX2_Vreftrim;
input		SP2HP_xTX2_activepkEn;
input		SP2HP_xTX2_busdivSel;
input		SP2HP_xTX2_chico_cksel;
input		SP2HP_xTX2_chico_pwrdnB;
input	[2:0]	SP2HP_xTX2_ctune;
input	[1:0]	SP2HP_xTX2_dccbiastrim;
input	[1:0]	SP2HP_xTX2_dccerrtrim;
input		SP2HP_xTX2_dccfix;
input	[2:0]	SP2HP_xTX2_gmtune;
input		SP2HP_xTX2_ovsdivEn;
input	[1:0]	SP2HP_xTX2_pdivSel;
input		SP2HP_xTX2_pwrdnB;
input		SP2HP_xTX2_selFourFive;
input		SP2HP_xTX2_sendidle;
input		SP2HP_xTX2_syncTxToUsrclk;
input		SP2HP_xTX2_tdccEn;
input		SP2HP_xTX2_tdccovrd;
input		SP2HP_xTX1_ACCCLK_ROTATEH;
input		SP2HP_xTX1_ACC_DIN_SEL;
input	[1:0]	SP2HP_xTX1_ACC_NSEL;
input	[7:0]	SP2HP_xTX1_ACC_OVERRIDE;
input		SP2HP_xTX1_ACC_OVERRIDE_EN;
input		SP2HP_xTX1_ACC_ROTATE;
input		SP2HP_xTX1_ACC_UPDNSW;
input		SP2HP_xTX1_Clk_pwrdnB;
input	[2:0]	SP2HP_xTX1_DrvPostCursor;
input	[2:0]	SP2HP_xTX1_DrvPreCursor;
input		SP2HP_xTX1_Drv_pwrdnB;
input	[2:0]	SP2HP_xTX1_Drvbiastrim;
input	[3:0]	SP2HP_xTX1_Drvswing;
input	[2:0]	SP2HP_xTX1_PI_captrim;
input		SP2HP_xTX1_PI_pwrdnB;
input	[1:0]	SP2HP_xTX1_PIbiasTrim;
input		SP2HP_xTX1_Resl_En;
input		SP2HP_xTX1_SSC_EN;
input	[8:0]	SP2HP_xTX1_SSC_OVERRIDE;
input		SP2HP_xTX1_SSC_OVERRIDE_EN;
input	[4:0]	SP2HP_xTX1_SSC_TSEL;
input		SP2HP_xTX1_Ser_pwrdnB;
input	[2:0]	SP2HP_xTX1_Serbiastrim;
input	[3:0]	SP2HP_xTX1_Vreftrim;
input		SP2HP_xTX1_activepkEn;
input		SP2HP_xTX1_busdivSel;
input		SP2HP_xTX1_chico_cksel;
input		SP2HP_xTX1_chico_pwrdnB;
input	[2:0]	SP2HP_xTX1_ctune;
input	[1:0]	SP2HP_xTX1_dccbiastrim;
input	[1:0]	SP2HP_xTX1_dccerrtrim;
input		SP2HP_xTX1_dccfix;
input	[2:0]	SP2HP_xTX1_gmtune;
input		SP2HP_xTX1_ovsdivEn;
input	[1:0]	SP2HP_xTX1_pdivSel;
input		SP2HP_xTX1_pwrdnB;
input		SP2HP_xTX1_selFourFive;
input		SP2HP_xTX1_sendidle;
input		SP2HP_xTX1_syncTxToUsrclk;
input		SP2HP_xTX1_tdccEn;
input		SP2HP_xTX1_tdccovrd;
input		SP2HP_xTX0_ACCCLK_ROTATEH;
input		SP2HP_xTX0_ACC_DIN_SEL;
input	[1:0]	SP2HP_xTX0_ACC_NSEL;
input	[7:0]	SP2HP_xTX0_ACC_OVERRIDE;
input		SP2HP_xTX0_ACC_OVERRIDE_EN;
input		SP2HP_xTX0_ACC_ROTATE;
input		SP2HP_xTX0_ACC_UPDNSW;
input		SP2HP_xTX0_Clk_pwrdnB;
input	[2:0]	SP2HP_xTX0_DrvPostCursor;
input	[2:0]	SP2HP_xTX0_DrvPreCursor;
input		SP2HP_xTX0_Drv_pwrdnB;
input	[2:0]	SP2HP_xTX0_Drvbiastrim;
input	[3:0]	SP2HP_xTX0_Drvswing;
input	[2:0]	SP2HP_xTX0_PI_captrim;
input		SP2HP_xTX0_PI_pwrdnB;
input	[1:0]	SP2HP_xTX0_PIbiasTrim;
input		SP2HP_xTX0_Resl_En;
input		SP2HP_xTX0_SSC_EN;
input	[8:0]	SP2HP_xTX0_SSC_OVERRIDE;
input		SP2HP_xTX0_SSC_OVERRIDE_EN;
input	[4:0]	SP2HP_xTX0_SSC_TSEL;
input		SP2HP_xTX0_Ser_pwrdnB;
input	[2:0]	SP2HP_xTX0_Serbiastrim;
input	[3:0]	SP2HP_xTX0_Vreftrim;
input		SP2HP_xTX0_activepkEn;
input		SP2HP_xTX0_busdivSel;
input		SP2HP_xTX0_chico_cksel;
input		SP2HP_xTX0_chico_pwrdnB;
input	[2:0]	SP2HP_xTX0_ctune;
input	[1:0]	SP2HP_xTX0_dccbiastrim;
input	[1:0]	SP2HP_xTX0_dccerrtrim;
input		SP2HP_xTX0_dccfix;
input	[2:0]	SP2HP_xTX0_gmtune;
input		SP2HP_xTX0_ovsdivEn;
input	[1:0]	SP2HP_xTX0_pdivSel;
input		SP2HP_xTX0_pwrdnB;
input		SP2HP_xTX0_selFourFive;
input		SP2HP_xTX0_sendidle;
input		SP2HP_xTX0_syncTxToUsrclk;
input		SP2HP_xTX0_tdccEn;
input		SP2HP_xTX0_tdccovrd;
input		SP2HP_xTX_SSC_Align;
input		clk_p;
input		fp2HP_L3RxBufClr;
input		fp2HP_L3RxCALSlide;
input		fp2HP_L3RxGearboxSlip;
input		fp2HP_L3RxPRBSCntClr;
input	[2:0]	fp2HP_L3RxPRBSTst;
input		fp2HP_L3RxPRBSZCntClr;
input		fp2HP_L3RxPolarity;
input		fp2HP_L3TxBitReverse;
input		fp2HP_L3TxBufClr;
input	[1:0]	fp2HP_L3TxDMux;
input		fp2HP_L3TxElecIdleAdj;
input	[1:0]	fp2HP_L3TxFlMux;
input		fp2HP_L3TxPCIEDetectRx;
input		fp2HP_L3TxPCIEElecIdle;
input	[2:0]	fp2HP_L3TxPMux;
input		fp2HP_L3TxPRBSErrCont;
input		fp2HP_L3TxPRBSErrOne;
input	[2:0]	fp2HP_L3TxPRBSTst;
input		fp2HP_L3TxPolarity;
input		fp2HP_L3TxSATAOOBComRESET;
input		fp2HP_L3TxSATAOOBComSAS;
input		fp2HP_L3TxSATAOOBComWAKE;
input	[7:0]	fp2HP_L3TxUsr8B10BDataK;
input	[7:0]	fp2HP_L3TxUsr8B10BDispMode;
input	[7:0]	fp2HP_L3TxUsr8B10BDispVal;
input	[79:0]	fp2HP_L3TxUsrData;
input	[2:0]	fp2HP_L3TxUsrGBHeader;
input	[6:0]	fp2HP_L3TxUsrGBSequence;
input		fp2HP_L3TxUsrGBStartSeq;
input		fp2HP_L2RxBufClr;
input		fp2HP_L2RxCALSlide;
input		fp2HP_L2RxGearboxSlip;
input		fp2HP_L2RxPRBSCntClr;
input	[2:0]	fp2HP_L2RxPRBSTst;
input		fp2HP_L2RxPRBSZCntClr;
input		fp2HP_L2RxPolarity;
input		fp2HP_L2TxBitReverse;
input		fp2HP_L2TxBufClr;
input	[1:0]	fp2HP_L2TxDMux;
input		fp2HP_L2TxElecIdleAdj;
input	[1:0]	fp2HP_L2TxFlMux;
input		fp2HP_L2TxPCIEDetectRx;
input		fp2HP_L2TxPCIEElecIdle;
input	[2:0]	fp2HP_L2TxPMux;
input		fp2HP_L2TxPRBSErrCont;
input		fp2HP_L2TxPRBSErrOne;
input	[2:0]	fp2HP_L2TxPRBSTst;
input		fp2HP_L2TxPolarity;
input		fp2HP_L2TxSATAOOBComRESET;
input		fp2HP_L2TxSATAOOBComSAS;
input		fp2HP_L2TxSATAOOBComWAKE;
input	[7:0]	fp2HP_L2TxUsr8B10BDataK;
input	[7:0]	fp2HP_L2TxUsr8B10BDispMode;
input	[7:0]	fp2HP_L2TxUsr8B10BDispVal;
input	[79:0]	fp2HP_L2TxUsrData;
input	[2:0]	fp2HP_L2TxUsrGBHeader;
input	[6:0]	fp2HP_L2TxUsrGBSequence;
input		fp2HP_L2TxUsrGBStartSeq;
input		fp2HP_L1RxBufClr;
input		fp2HP_L1RxCALSlide;
input		fp2HP_L1RxGearboxSlip;
input		fp2HP_L1RxPRBSCntClr;
input	[2:0]	fp2HP_L1RxPRBSTst;
input		fp2HP_L1RxPRBSZCntClr;
input		fp2HP_L1RxPolarity;
input		fp2HP_L1TxBitReverse;
input		fp2HP_L1TxBufClr;
input	[1:0]	fp2HP_L1TxDMux;
input		fp2HP_L1TxElecIdleAdj;
input	[1:0]	fp2HP_L1TxFlMux;
input		fp2HP_L1TxPCIEDetectRx;
input		fp2HP_L1TxPCIEElecIdle;
input	[2:0]	fp2HP_L1TxPMux;
input		fp2HP_L1TxPRBSErrCont;
input		fp2HP_L1TxPRBSErrOne;
input	[2:0]	fp2HP_L1TxPRBSTst;
input		fp2HP_L1TxPolarity;
input		fp2HP_L1TxSATAOOBComRESET;
input		fp2HP_L1TxSATAOOBComSAS;
input		fp2HP_L1TxSATAOOBComWAKE;
input	[7:0]	fp2HP_L1TxUsr8B10BDataK;
input	[7:0]	fp2HP_L1TxUsr8B10BDispMode;
input	[7:0]	fp2HP_L1TxUsr8B10BDispVal;
input	[79:0]	fp2HP_L1TxUsrData;
input	[2:0]	fp2HP_L1TxUsrGBHeader;
input	[6:0]	fp2HP_L1TxUsrGBSequence;
input		fp2HP_L1TxUsrGBStartSeq;
input		fp2HP_L0RxBufClr;
input		fp2HP_L0RxCALSlide;
input		fp2HP_L0RxGearboxSlip;
input		fp2HP_L0RxPRBSCntClr;
input	[2:0]	fp2HP_L0RxPRBSTst;
input		fp2HP_L0RxPRBSZCntClr;
input		fp2HP_L0RxPolarity;
input		fp2HP_L0TxBitReverse;
input		fp2HP_L0TxBufClr;
input	[1:0]	fp2HP_L0TxDMux;
input		fp2HP_L0TxElecIdleAdj;
input	[1:0]	fp2HP_L0TxFlMux;
input		fp2HP_L0TxPCIEDetectRx;
input		fp2HP_L0TxPCIEElecIdle;
input	[2:0]	fp2HP_L0TxPMux;
input		fp2HP_L0TxPRBSErrCont;
input		fp2HP_L0TxPRBSErrOne;
input	[2:0]	fp2HP_L0TxPRBSTst;
input		fp2HP_L0TxPolarity;
input		fp2HP_L0TxSATAOOBComRESET;
input		fp2HP_L0TxSATAOOBComSAS;
input		fp2HP_L0TxSATAOOBComWAKE;
input	[7:0]	fp2HP_L0TxUsr8B10BDataK;
input	[7:0]	fp2HP_L0TxUsr8B10BDispMode;
input	[7:0]	fp2HP_L0TxUsr8B10BDispVal;
input	[79:0]	fp2HP_L0TxUsrData;
input	[2:0]	fp2HP_L0TxUsrGBHeader;
input	[6:0]	fp2HP_L0TxUsrGBSequence;
input		fp2HP_L0TxUsrGBStartSeq;
input		fp2HP_UsrRst_N;
input		fp2HP_UsrRxRst_N;
input		fp2HP_UsrTxRst_N;
input		fp2HP_pcs_usr_resetB;
input	[31:0]	pbus_addr;
input		pbus_req;
input	[31:0]	pbus_wdata;
input		pbus_write;
input		rst_p_n;
input		xCMU_grefclk;

parameter  cfg_wrdly = 2'b0;
parameter serdes_iso_en = 1'b0;
parameter cfg_mux_fp_pcie_L3 = 1'b0;
parameter cfg_mux_fp_pcie_L2 = 1'b0;
parameter cfg_mux_fp_pcie_L1 = 1'b0;
parameter cfg_mux_fp_pcie_L0 = 1'b0;
parameter cfg_serdes_dbgck_sel = 1'b0;
parameter cfg_serdes_by_reg = 1'b0;
parameter cfg_mux_fp_pcie_common = 1'b0;

// PCS CFG Common Registers, Offset = 15'h4000
parameter SYSTEMRESET                 = 16'h0001;    // Offset = 15'h4000 Attributes : RW   
parameter MODESET                     = 16'h0007;    // Offset = 15'h4001 Attributes : RW   
parameter RXLDUNIFORMCLKSEL           = 16'h0000;    // Offset = 15'h4002 Attributes : RW   
parameter RXLDSTATUS                  = 16'h0000;    // Offset = 15'h4003 Attributes : RO   
parameter LANEEN                      = 16'h000f;    // Offset = 15'h4004 Attributes : RW   
parameter SSCENX4                     = 16'h0000;    // Offset = 15'h4005 Attributes : RW   
parameter SOFTRST                     = 16'h0000;    // Offset = 15'h4008 Attributes : RW   
parameter TXDETRX1                    = 16'h0048;    // Offset = 15'h4010 Attributes : RW   
parameter TXDETRX2                    = 16'h00a2;    // Offset = 15'h4011 Attributes : RW   
parameter PININITT                    = 16'd2000;    // Offset = 15'h4020 Attributes : RW   
parameter PONPWRINTVALT               = 16'd2000;    // Offset = 15'h4021 Attributes : RW   
parameter PONPRERESCALT               = 16'd2000;    // Offset = 15'h4022 Attributes : RW   
parameter PONRESCALHIT                = 16'd1000;    // Offset = 15'h4023 Attributes : RW   
parameter PONRESCALLOT                = 16'd0200;    // Offset = 15'h4024 Attributes : RW   
parameter PONPREPLLDETT               = 16'd1000;    // Offset = 15'h4025 Attributes : RW   
parameter PONPLLDETT                  = 16'd3000;    // Offset = 15'h4026 Attributes : RW   
parameter PONCHGCLKT1                 = 16'h0fff;    // Offset = 15'h4027 Attributes : RW   
parameter PONCHGCLKT2                 = 16'd3000;    // Offset = 15'h4028 Attributes : RW   
parameter PONOFSTCALHIT               = 16'd1000;    // Offset = 15'h4029 Attributes : RW   
parameter POWERONCTRL                 = 16'h0000;    // Offset = 15'h402E Attributes : RW   
parameter POWERONSTATUS               = 16'h0000;    // Offset = 15'h402F Attributes : RO   
parameter PONOFSTCALLOT               = 16'd0200;    // Offset = 15'h402a Attributes : RW   
parameter PONPREDFECALT               = 16'd2000;    // Offset = 15'h402b Attributes : RW   
parameter PONDFECALT                  = 16'd1000;    // Offset = 15'h402c Attributes : RW   
parameter RESCALCTRL                  = 16'h0000;    // Offset = 15'h4030 Attributes : RW   
parameter RESCALSTATUS                = 16'h0000;    // Offset = 15'h4031 Attributes : RO   
parameter TxPhaseAlignT               = 16'd8000;    // Offset = 15'h4040 Attributes : RW   
parameter PIPECTRL                    = 16'h0000;    // Offset = 15'h4050 Attributes : RW   
parameter PIPERATESET                 = 16'h0000;    // Offset = 15'h4051 Attributes : RO   

// PCS CFG Lane Registers, Offset = 15'h0000(Lane0) 15'h0200(Lane1) 15'h0400(Lane2) 15'h0600(Lane3) 15'h1000(Broadcast)
parameter L0_TXDMUX                   = 16'h0101;    // Offset = 15'h000 Attributes : RW   
parameter L0_TXOOBSET                 = 16'h1561;    // Offset = 15'h001 Attributes : RW   
parameter L0_TXOOBSEND                = 16'h0000;    // Offset = 15'h002 Attributes : WST   
parameter L0_TXOOBSENDSTATUS          = 16'h0000;    // Offset = 15'h003 Attributes : RO   
parameter L0_TXPHASET                 = 16'h0003;    // Offset = 15'h004 Attributes : RW   
parameter L0_TXPHACLR                 = 16'h0000;    // Offset = 15'h005 Attributes : RW   
parameter L0_TXPHASTATUS              = 16'h0000;    // Offset = 15'h006 Attributes : RO   
parameter L0_TXPMUX                   = 16'h0002;    // Offset = 15'h008 Attributes : RW   
parameter L0_TXPRBSGENSET             = 16'h0001;    // Offset = 15'h00C Attributes : RW   
parameter L0_TXPRBSGENDEBUG           = 16'h0000;    // Offset = 15'h00D Attributes : RW   
parameter L0_TXPRBSGENPATTEN1         = 16'h03ff;    // Offset = 15'h010 Attributes : RW   
parameter L0_TXPRBSGENPATTEN2         = 16'h03ff;    // Offset = 15'h011 Attributes : RW   
parameter L0_TXPRBSGENPATTEN3         = 16'h0000;    // Offset = 15'h012 Attributes : RW   
parameter L0_TXPRBSGENPATTEN4         = 16'h0000;    // Offset = 15'h013 Attributes : RW   
parameter L0_TXENC8TO10               = 16'h0001;    // Offset = 15'h014 Attributes : RW   
parameter L0_TXENC8TO10DISP           = 16'h0000;    // Offset = 15'h015 Attributes : RO   
parameter L0_TXENC8TO10ERRCNT         = 16'h0000;    // Offset = 15'h016 Attributes : RO   
parameter L0_TXENC8TO10ERRCNTCLR      = 16'h0000;    // Offset = 15'h017 Attributes : RW   
parameter L0_TXGEARBOX                = 16'h0000;    // Offset = 15'h018 Attributes : RW   
parameter L0_TXENC4TO5                = 16'h0000;    // Offset = 15'h019 Attributes : RW   
parameter L0_TXFLMUX                  = 16'h0001;    // Offset = 15'h01C Attributes : RW   
parameter L0_TXUIA                    = 16'h0000;    // Offset = 15'h020 Attributes : RW   
parameter L0_RXOVRSMPLSET             = 16'h2002;    // Offset = 15'h100 Attributes : RW   
parameter L0_RXOVRSMPLERRCNT          = 16'h0000;    // Offset = 15'h101 Attributes : RO   
parameter L0_RXOVRSMPLERRCNTCLR       = 16'h0000;    // Offset = 15'h102 Attributes : RW   
parameter L0_RXOOBBURST               = 16'h0603;    // Offset = 15'h104 Attributes : RW   
parameter L0_RXOOBCOMINIT             = 16'h2208;    // Offset = 15'h105 Attributes : RW   
parameter L0_RXOOBCOMSAS              = 16'h7525;    // Offset = 15'h106 Attributes : RW   
parameter L0_RXOOBCOMWAKE             = 16'h0603;    // Offset = 15'h107 Attributes : RW   
parameter L0_RXOOBSET                 = 16'h0006;    // Offset = 15'h108 Attributes : RW   
parameter L0_RXOOBSTATUS              = 16'h0000;    // Offset = 15'h109 Attributes : RO   
parameter L0_RXOOBCOMINITCNT          = 16'h0000;    // Offset = 15'h10A Attributes : RO   
parameter L0_RXOOBCOMSASCNT           = 16'h0000;    // Offset = 15'h10B Attributes : RO   
parameter L0_RXOOBCOMWAKECNT          = 16'h0000;    // Offset = 15'h10C Attributes : RO   
parameter L0_RXOOBCNTCLR              = 16'h0000;    // Offset = 15'h10D Attributes : RW   
parameter L0_RXPRBSCHK                = 16'h0001;    // Offset = 15'h110 Attributes : RW   
parameter L0_RXPRBSCHKERRCNT          = 16'h0000;    // Offset = 15'h111 Attributes : RO   
parameter L0_RXPRBSZEROCNT            = 16'h0000;    // Offset = 15'h112 Attributes : RO   
parameter L0_RXPRBSCHKCNTCLR          = 16'h0000;    // Offset = 15'h113 Attributes : RW   
parameter L0_RXPRBSCHKPATTEN1         = 16'h03ff;    // Offset = 15'h114 Attributes : RW   
parameter L0_RXPRBSCHKPATTEN2         = 16'h03ff;    // Offset = 15'h115 Attributes : RW   
parameter L0_RXPRBSCHKPATTEN3         = 16'h0000;    // Offset = 15'h116 Attributes : RW   
parameter L0_RXPRBSCHKPATTEN4         = 16'h0000;    // Offset = 15'h117 Attributes : RW   
parameter L0_RX8B10BCAD               = 16'hc3ff;    // Offset = 15'h120 Attributes : RW   
parameter L0_RX8B10BCADMCOMMA         = 16'h2283;    // Offset = 15'h121 Attributes : RW   
parameter L0_RX8B10BCADPCOMMA         = 16'h217c;    // Offset = 15'h122 Attributes : RW   
parameter L0_RX8B10BCADSLIDE          = 16'h0000;    // Offset = 15'h123 Attributes : RW   
parameter L0_RX8B10BDEC               = 16'h0001;    // Offset = 15'h124 Attributes : RW   
parameter L0_RX8B10BDECCOMMA          = 16'h0000;    // Offset = 15'h125 Attributes : RW   
parameter L0_RX8B10BSYNC              = 16'h5111;    // Offset = 15'h128 Attributes : RW   
parameter L0_RX8B10BSTATUS            = 16'h0000;    // Offset = 15'h129 Attributes : RO   
parameter L0_RX4B5BSET                = 16'h0000;    // Offset = 15'h12B Attributes : RW   
parameter L0_RX4B5BSD                 = 16'h0223;    // Offset = 15'h12C Attributes : RW   
parameter L0_RX4B5BED                 = 16'h0396;    // Offset = 15'h12D Attributes : RW   
parameter L0_RXPMUX                   = 16'h0001;    // Offset = 15'h12F Attributes : RW   
parameter L0_RXLDBUF                  = 16'h0000;    // Offset = 15'h130 Attributes : RW   
parameter L0_RXLDBUFSEQ1              = 16'h0000;    // Offset = 15'h131 Attributes : RW   
parameter L0_RXLDBUFSEQ2              = 16'h0000;    // Offset = 15'h132 Attributes : RW   
parameter L0_RXLDBUFSEQ3              = 16'h0000;    // Offset = 15'h133 Attributes : RW   
parameter L0_RXLDBUFSEQ4              = 16'h0000;    // Offset = 15'h134 Attributes : RW   
parameter L0_RXLDBUFSEQEN             = 16'hf1ff;    // Offset = 15'h135 Attributes : RW   
parameter L0_RXEBUF                   = 16'h0001;    // Offset = 15'h138 Attributes : RW   
parameter L0_RXEBUFCLR                = 16'h0000;    // Offset = 15'h139 Attributes : RW   
parameter L0_RXCLKCOR                 = 16'h0101;    // Offset = 15'h13A Attributes : RW   
parameter L0_RXCLKCORSEQ1             = 16'h011c;    // Offset = 15'h13C Attributes : RW   
parameter L0_RXCLKCORSEQ2             = 16'h0000;    // Offset = 15'h13D Attributes : RW   
parameter L0_RXCLKCORSEQ3             = 16'h0000;    // Offset = 15'h13E Attributes : RW   
parameter L0_RXCLKCORSEQ4             = 16'h0000;    // Offset = 15'h13F Attributes : RW   
parameter L0_RXGEARBOX                = 16'h0000;    // Offset = 15'h140 Attributes : RW   
parameter L0_RXGEARBOXSLIP            = 16'h0000;    // Offset = 15'h141 Attributes : RW   
parameter L0_RXGEARBOXSTATUS          = 16'h0000;    // Offset = 15'h142 Attributes : RO   
parameter L0_RXUIA                    = 16'h0000;    // Offset = 15'h144 Attributes : RW   
parameter L0_PCSCMU                   = 16'hd812;    // Offset = 15'h148 Attributes : RW   
parameter L0_PMAUBRDSET               = 16'h0000;    // Offset = 15'h151 Attributes : RW   
parameter L0_PMAUBRDRSLT              = 16'h0000;    // Offset = 15'h152 Attributes : RO   
parameter L0_PMAUBOFCALSET            = 16'h0000;    // Offset = 15'h153 Attributes : RW   
parameter L0_PMAUBOFCALRSLT           = 16'h0000;    // Offset = 15'h154 Attributes : RO   
parameter L0_PMAUBPHASET              = 16'h0000;    // Offset = 15'h155 Attributes : RW   
parameter L0_PMAUBPHARSLT             = 16'h0000;    // Offset = 15'h156 Attributes : RO   
parameter L0_PCSRMUSRST               = 16'h0000;    // Offset = 15'h158 Attributes : RW   

parameter L1_TXDMUX                   = 16'h0101;    // Offset = 15'h200 Attributes : RW   
parameter L1_TXOOBSET                 = 16'h1561;    // Offset = 15'h201 Attributes : RW   
parameter L1_TXOOBSEND                = 16'h0000;    // Offset = 15'h202 Attributes : WST   
parameter L1_TXOOBSENDSTATUS          = 16'h0000;    // Offset = 15'h203 Attributes : RO   
parameter L1_TXPHASET                 = 16'h0003;    // Offset = 15'h204 Attributes : RW   
parameter L1_TXPHACLR                 = 16'h0000;    // Offset = 15'h205 Attributes : RW   
parameter L1_TXPHASTATUS              = 16'h0000;    // Offset = 15'h206 Attributes : RO   
parameter L1_TXPMUX                   = 16'h0002;    // Offset = 15'h208 Attributes : RW   
parameter L1_TXPRBSGENSET             = 16'h0001;    // Offset = 15'h20C Attributes : RW   
parameter L1_TXPRBSGENDEBUG           = 16'h0000;    // Offset = 15'h20D Attributes : RW   
parameter L1_TXPRBSGENPATTEN1         = 16'h03ff;    // Offset = 15'h210 Attributes : RW   
parameter L1_TXPRBSGENPATTEN2         = 16'h03ff;    // Offset = 15'h211 Attributes : RW   
parameter L1_TXPRBSGENPATTEN3         = 16'h0000;    // Offset = 15'h212 Attributes : RW   
parameter L1_TXPRBSGENPATTEN4         = 16'h0000;    // Offset = 15'h213 Attributes : RW   
parameter L1_TXENC8TO10               = 16'h0001;    // Offset = 15'h214 Attributes : RW   
parameter L1_TXENC8TO10DISP           = 16'h0000;    // Offset = 15'h215 Attributes : RO   
parameter L1_TXENC8TO10ERRCNT         = 16'h0000;    // Offset = 15'h216 Attributes : RO   
parameter L1_TXENC8TO10ERRCNTCLR      = 16'h0000;    // Offset = 15'h217 Attributes : RW   
parameter L1_TXGEARBOX                = 16'h0000;    // Offset = 15'h218 Attributes : RW   
parameter L1_TXENC4TO5                = 16'h0000;    // Offset = 15'h219 Attributes : RW   
parameter L1_TXFLMUX                  = 16'h0001;    // Offset = 15'h21C Attributes : RW   
parameter L1_TXUIA                    = 16'h0000;    // Offset = 15'h220 Attributes : RW   
parameter L1_RXOVRSMPLSET             = 16'h2002;    // Offset = 15'h300 Attributes : RW   
parameter L1_RXOVRSMPLERRCNT          = 16'h0000;    // Offset = 15'h301 Attributes : RO   
parameter L1_RXOVRSMPLERRCNTCLR       = 16'h0000;    // Offset = 15'h302 Attributes : RW   
parameter L1_RXOOBBURST               = 16'h0603;    // Offset = 15'h304 Attributes : RW   
parameter L1_RXOOBCOMINIT             = 16'h2208;    // Offset = 15'h305 Attributes : RW   
parameter L1_RXOOBCOMSAS              = 16'h7525;    // Offset = 15'h306 Attributes : RW   
parameter L1_RXOOBCOMWAKE             = 16'h0603;    // Offset = 15'h307 Attributes : RW   
parameter L1_RXOOBSET                 = 16'h0006;    // Offset = 15'h308 Attributes : RW   
parameter L1_RXOOBSTATUS              = 16'h0000;    // Offset = 15'h309 Attributes : RO   
parameter L1_RXOOBCOMINITCNT          = 16'h0000;    // Offset = 15'h30A Attributes : RO   
parameter L1_RXOOBCOMSASCNT           = 16'h0000;    // Offset = 15'h30B Attributes : RO   
parameter L1_RXOOBCOMWAKECNT          = 16'h0000;    // Offset = 15'h30C Attributes : RO   
parameter L1_RXOOBCNTCLR              = 16'h0000;    // Offset = 15'h30D Attributes : RW   
parameter L1_RXPRBSCHK                = 16'h0001;    // Offset = 15'h310 Attributes : RW   
parameter L1_RXPRBSCHKERRCNT          = 16'h0000;    // Offset = 15'h311 Attributes : RO   
parameter L1_RXPRBSZEROCNT            = 16'h0000;    // Offset = 15'h312 Attributes : RO   
parameter L1_RXPRBSCHKCNTCLR          = 16'h0000;    // Offset = 15'h313 Attributes : RW   
parameter L1_RXPRBSCHKPATTEN1         = 16'h03ff;    // Offset = 15'h314 Attributes : RW   
parameter L1_RXPRBSCHKPATTEN2         = 16'h03ff;    // Offset = 15'h315 Attributes : RW   
parameter L1_RXPRBSCHKPATTEN3         = 16'h0000;    // Offset = 15'h316 Attributes : RW   
parameter L1_RXPRBSCHKPATTEN4         = 16'h0000;    // Offset = 15'h317 Attributes : RW   
parameter L1_RX8B10BCAD               = 16'hc3ff;    // Offset = 15'h320 Attributes : RW   
parameter L1_RX8B10BCADMCOMMA         = 16'h2283;    // Offset = 15'h321 Attributes : RW   
parameter L1_RX8B10BCADPCOMMA         = 16'h217c;    // Offset = 15'h322 Attributes : RW   
parameter L1_RX8B10BCADSLIDE          = 16'h0000;    // Offset = 15'h323 Attributes : RW   
parameter L1_RX8B10BDEC               = 16'h0001;    // Offset = 15'h324 Attributes : RW   
parameter L1_RX8B10BDECCOMMA          = 16'h0000;    // Offset = 15'h325 Attributes : RW   
parameter L1_RX8B10BSYNC              = 16'h5111;    // Offset = 15'h328 Attributes : RW   
parameter L1_RX8B10BSTATUS            = 16'h0000;    // Offset = 15'h329 Attributes : RO   
parameter L1_RX4B5BSET                = 16'h0000;    // Offset = 15'h32B Attributes : RW   
parameter L1_RX4B5BSD                 = 16'h0223;    // Offset = 15'h32C Attributes : RW   
parameter L1_RX4B5BED                 = 16'h0396;    // Offset = 15'h32D Attributes : RW   
parameter L1_RXPMUX                   = 16'h0001;    // Offset = 15'h32F Attributes : RW   
parameter L1_RXLDBUF                  = 16'h0000;    // Offset = 15'h330 Attributes : RW   
parameter L1_RXLDBUFSEQ1              = 16'h0000;    // Offset = 15'h331 Attributes : RW   
parameter L1_RXLDBUFSEQ2              = 16'h0000;    // Offset = 15'h332 Attributes : RW   
parameter L1_RXLDBUFSEQ3              = 16'h0000;    // Offset = 15'h333 Attributes : RW   
parameter L1_RXLDBUFSEQ4              = 16'h0000;    // Offset = 15'h334 Attributes : RW   
parameter L1_RXLDBUFSEQEN             = 16'hf1ff;    // Offset = 15'h335 Attributes : RW   
parameter L1_RXEBUF                   = 16'h0001;    // Offset = 15'h338 Attributes : RW   
parameter L1_RXEBUFCLR                = 16'h0000;    // Offset = 15'h339 Attributes : RW   
parameter L1_RXCLKCOR                 = 16'h0101;    // Offset = 15'h33A Attributes : RW   
parameter L1_RXCLKCORSEQ1             = 16'h011c;    // Offset = 15'h33C Attributes : RW   
parameter L1_RXCLKCORSEQ2             = 16'h0000;    // Offset = 15'h33D Attributes : RW   
parameter L1_RXCLKCORSEQ3             = 16'h0000;    // Offset = 15'h33E Attributes : RW   
parameter L1_RXCLKCORSEQ4             = 16'h0000;    // Offset = 15'h33F Attributes : RW   
parameter L1_RXGEARBOX                = 16'h0000;    // Offset = 15'h340 Attributes : RW   
parameter L1_RXGEARBOXSLIP            = 16'h0000;    // Offset = 15'h341 Attributes : RW   
parameter L1_RXGEARBOXSTATUS          = 16'h0000;    // Offset = 15'h342 Attributes : RO   
parameter L1_RXUIA                    = 16'h0000;    // Offset = 15'h344 Attributes : RW   
parameter L1_PCSCMU                   = 16'hd812;    // Offset = 15'h348 Attributes : RW   
parameter L1_PMAUBRDSET               = 16'h0000;    // Offset = 15'h351 Attributes : RW   
parameter L1_PMAUBRDRSLT              = 16'h0000;    // Offset = 15'h352 Attributes : RO   
parameter L1_PMAUBOFCALSET            = 16'h0000;    // Offset = 15'h353 Attributes : RW   
parameter L1_PMAUBOFCALRSLT           = 16'h0000;    // Offset = 15'h354 Attributes : RO   
parameter L1_PMAUBPHASET              = 16'h0000;    // Offset = 15'h355 Attributes : RW   
parameter L1_PMAUBPHARSLT             = 16'h0000;    // Offset = 15'h356 Attributes : RO   
parameter L1_PCSRMUSRST               = 16'h0000;    // Offset = 15'h358 Attributes : RW   

parameter L2_TXDMUX                   = 16'h0101;    // Offset = 15'h400 Attributes : RW   
parameter L2_TXOOBSET                 = 16'h1561;    // Offset = 15'h401 Attributes : RW   
parameter L2_TXOOBSEND                = 16'h0000;    // Offset = 15'h402 Attributes : WST   
parameter L2_TXOOBSENDSTATUS          = 16'h0000;    // Offset = 15'h403 Attributes : RO   
parameter L2_TXPHASET                 = 16'h0003;    // Offset = 15'h404 Attributes : RW   
parameter L2_TXPHACLR                 = 16'h0000;    // Offset = 15'h405 Attributes : RW   
parameter L2_TXPHASTATUS              = 16'h0000;    // Offset = 15'h406 Attributes : RO   
parameter L2_TXPMUX                   = 16'h0002;    // Offset = 15'h408 Attributes : RW   
parameter L2_TXPRBSGENSET             = 16'h0001;    // Offset = 15'h40C Attributes : RW   
parameter L2_TXPRBSGENDEBUG           = 16'h0000;    // Offset = 15'h40D Attributes : RW   
parameter L2_TXPRBSGENPATTEN1         = 16'h03ff;    // Offset = 15'h410 Attributes : RW   
parameter L2_TXPRBSGENPATTEN2         = 16'h03ff;    // Offset = 15'h411 Attributes : RW   
parameter L2_TXPRBSGENPATTEN3         = 16'h0000;    // Offset = 15'h412 Attributes : RW   
parameter L2_TXPRBSGENPATTEN4         = 16'h0000;    // Offset = 15'h413 Attributes : RW   
parameter L2_TXENC8TO10               = 16'h0001;    // Offset = 15'h414 Attributes : RW   
parameter L2_TXENC8TO10DISP           = 16'h0000;    // Offset = 15'h415 Attributes : RO   
parameter L2_TXENC8TO10ERRCNT         = 16'h0000;    // Offset = 15'h416 Attributes : RO   
parameter L2_TXENC8TO10ERRCNTCLR      = 16'h0000;    // Offset = 15'h417 Attributes : RW   
parameter L2_TXGEARBOX                = 16'h0000;    // Offset = 15'h418 Attributes : RW   
parameter L2_TXENC4TO5                = 16'h0000;    // Offset = 15'h419 Attributes : RW   
parameter L2_TXFLMUX                  = 16'h0001;    // Offset = 15'h41C Attributes : RW   
parameter L2_TXUIA                    = 16'h0000;    // Offset = 15'h420 Attributes : RW   
parameter L2_RXOVRSMPLSET             = 16'h2002;    // Offset = 15'h500 Attributes : RW   
parameter L2_RXOVRSMPLERRCNT          = 16'h0000;    // Offset = 15'h501 Attributes : RO   
parameter L2_RXOVRSMPLERRCNTCLR       = 16'h0000;    // Offset = 15'h502 Attributes : RW   
parameter L2_RXOOBBURST               = 16'h0603;    // Offset = 15'h504 Attributes : RW   
parameter L2_RXOOBCOMINIT             = 16'h2208;    // Offset = 15'h505 Attributes : RW   
parameter L2_RXOOBCOMSAS              = 16'h7525;    // Offset = 15'h506 Attributes : RW   
parameter L2_RXOOBCOMWAKE             = 16'h0603;    // Offset = 15'h507 Attributes : RW   
parameter L2_RXOOBSET                 = 16'h0006;    // Offset = 15'h508 Attributes : RW   
parameter L2_RXOOBSTATUS              = 16'h0000;    // Offset = 15'h509 Attributes : RO   
parameter L2_RXOOBCOMINITCNT          = 16'h0000;    // Offset = 15'h50A Attributes : RO   
parameter L2_RXOOBCOMSASCNT           = 16'h0000;    // Offset = 15'h50B Attributes : RO   
parameter L2_RXOOBCOMWAKECNT          = 16'h0000;    // Offset = 15'h50C Attributes : RO   
parameter L2_RXOOBCNTCLR              = 16'h0000;    // Offset = 15'h50D Attributes : RW   
parameter L2_RXPRBSCHK                = 16'h0001;    // Offset = 15'h510 Attributes : RW   
parameter L2_RXPRBSCHKERRCNT          = 16'h0000;    // Offset = 15'h511 Attributes : RO   
parameter L2_RXPRBSZEROCNT            = 16'h0000;    // Offset = 15'h512 Attributes : RO   
parameter L2_RXPRBSCHKCNTCLR          = 16'h0000;    // Offset = 15'h513 Attributes : RW   
parameter L2_RXPRBSCHKPATTEN1         = 16'h03ff;    // Offset = 15'h514 Attributes : RW   
parameter L2_RXPRBSCHKPATTEN2         = 16'h03ff;    // Offset = 15'h515 Attributes : RW   
parameter L2_RXPRBSCHKPATTEN3         = 16'h0000;    // Offset = 15'h516 Attributes : RW   
parameter L2_RXPRBSCHKPATTEN4         = 16'h0000;    // Offset = 15'h517 Attributes : RW   
parameter L2_RX8B10BCAD               = 16'hc3ff;    // Offset = 15'h520 Attributes : RW   
parameter L2_RX8B10BCADMCOMMA         = 16'h2283;    // Offset = 15'h521 Attributes : RW   
parameter L2_RX8B10BCADPCOMMA         = 16'h217c;    // Offset = 15'h522 Attributes : RW   
parameter L2_RX8B10BCADSLIDE          = 16'h0000;    // Offset = 15'h523 Attributes : RW   
parameter L2_RX8B10BDEC               = 16'h0001;    // Offset = 15'h524 Attributes : RW   
parameter L2_RX8B10BDECCOMMA          = 16'h0000;    // Offset = 15'h525 Attributes : RW   
parameter L2_RX8B10BSYNC              = 16'h5111;    // Offset = 15'h528 Attributes : RW   
parameter L2_RX8B10BSTATUS            = 16'h0000;    // Offset = 15'h529 Attributes : RO   
parameter L2_RX4B5BSET                = 16'h0000;    // Offset = 15'h52B Attributes : RW   
parameter L2_RX4B5BSD                 = 16'h0223;    // Offset = 15'h52C Attributes : RW   
parameter L2_RX4B5BED                 = 16'h0396;    // Offset = 15'h52D Attributes : RW   
parameter L2_RXPMUX                   = 16'h0001;    // Offset = 15'h52F Attributes : RW   
parameter L2_RXLDBUF                  = 16'h0000;    // Offset = 15'h530 Attributes : RW   
parameter L2_RXLDBUFSEQ1              = 16'h0000;    // Offset = 15'h531 Attributes : RW   
parameter L2_RXLDBUFSEQ2              = 16'h0000;    // Offset = 15'h532 Attributes : RW   
parameter L2_RXLDBUFSEQ3              = 16'h0000;    // Offset = 15'h533 Attributes : RW   
parameter L2_RXLDBUFSEQ4              = 16'h0000;    // Offset = 15'h534 Attributes : RW   
parameter L2_RXLDBUFSEQEN             = 16'hf1ff;    // Offset = 15'h535 Attributes : RW   
parameter L2_RXEBUF                   = 16'h0001;    // Offset = 15'h538 Attributes : RW   
parameter L2_RXEBUFCLR                = 16'h0000;    // Offset = 15'h539 Attributes : RW   
parameter L2_RXCLKCOR                 = 16'h0101;    // Offset = 15'h53A Attributes : RW   
parameter L2_RXCLKCORSEQ1             = 16'h011c;    // Offset = 15'h53C Attributes : RW   
parameter L2_RXCLKCORSEQ2             = 16'h0000;    // Offset = 15'h53D Attributes : RW   
parameter L2_RXCLKCORSEQ3             = 16'h0000;    // Offset = 15'h53E Attributes : RW   
parameter L2_RXCLKCORSEQ4             = 16'h0000;    // Offset = 15'h53F Attributes : RW   
parameter L2_RXGEARBOX                = 16'h0000;    // Offset = 15'h540 Attributes : RW   
parameter L2_RXGEARBOXSLIP            = 16'h0000;    // Offset = 15'h541 Attributes : RW   
parameter L2_RXGEARBOXSTATUS          = 16'h0000;    // Offset = 15'h542 Attributes : RO   
parameter L2_RXUIA                    = 16'h0000;    // Offset = 15'h544 Attributes : RW   
parameter L2_PCSCMU                   = 16'hd812;    // Offset = 15'h548 Attributes : RW   
parameter L2_PMAUBRDSET               = 16'h0000;    // Offset = 15'h551 Attributes : RW   
parameter L2_PMAUBRDRSLT              = 16'h0000;    // Offset = 15'h552 Attributes : RO   
parameter L2_PMAUBOFCALSET            = 16'h0000;    // Offset = 15'h553 Attributes : RW   
parameter L2_PMAUBOFCALRSLT           = 16'h0000;    // Offset = 15'h554 Attributes : RO   
parameter L2_PMAUBPHASET              = 16'h0000;    // Offset = 15'h555 Attributes : RW   
parameter L2_PMAUBPHARSLT             = 16'h0000;    // Offset = 15'h556 Attributes : RO   
parameter L2_PCSRMUSRST               = 16'h0000;    // Offset = 15'h558 Attributes : RW   

parameter L3_TXDMUX                   = 16'h0101;    // Offset = 15'h600 Attributes : RW   
parameter L3_TXOOBSET                 = 16'h1561;    // Offset = 15'h601 Attributes : RW   
parameter L3_TXOOBSEND                = 16'h0000;    // Offset = 15'h602 Attributes : WST   
parameter L3_TXOOBSENDSTATUS          = 16'h0000;    // Offset = 15'h603 Attributes : RO   
parameter L3_TXPHASET                 = 16'h0003;    // Offset = 15'h604 Attributes : RW   
parameter L3_TXPHACLR                 = 16'h0000;    // Offset = 15'h605 Attributes : RW   
parameter L3_TXPHASTATUS              = 16'h0000;    // Offset = 15'h606 Attributes : RO   
parameter L3_TXPMUX                   = 16'h0002;    // Offset = 15'h608 Attributes : RW   
parameter L3_TXPRBSGENSET             = 16'h0001;    // Offset = 15'h60C Attributes : RW   
parameter L3_TXPRBSGENDEBUG           = 16'h0000;    // Offset = 15'h60D Attributes : RW   
parameter L3_TXPRBSGENPATTEN1         = 16'h03ff;    // Offset = 15'h610 Attributes : RW   
parameter L3_TXPRBSGENPATTEN2         = 16'h03ff;    // Offset = 15'h611 Attributes : RW   
parameter L3_TXPRBSGENPATTEN3         = 16'h0000;    // Offset = 15'h612 Attributes : RW   
parameter L3_TXPRBSGENPATTEN4         = 16'h0000;    // Offset = 15'h613 Attributes : RW   
parameter L3_TXENC8TO10               = 16'h0001;    // Offset = 15'h614 Attributes : RW   
parameter L3_TXENC8TO10DISP           = 16'h0000;    // Offset = 15'h615 Attributes : RO   
parameter L3_TXENC8TO10ERRCNT         = 16'h0000;    // Offset = 15'h616 Attributes : RO   
parameter L3_TXENC8TO10ERRCNTCLR      = 16'h0000;    // Offset = 15'h617 Attributes : RW   
parameter L3_TXGEARBOX                = 16'h0000;    // Offset = 15'h618 Attributes : RW   
parameter L3_TXENC4TO5                = 16'h0000;    // Offset = 15'h619 Attributes : RW   
parameter L3_TXFLMUX                  = 16'h0001;    // Offset = 15'h61C Attributes : RW   
parameter L3_TXUIA                    = 16'h0000;    // Offset = 15'h620 Attributes : RW   
parameter L3_RXOVRSMPLSET             = 16'h2002;    // Offset = 15'h700 Attributes : RW   
parameter L3_RXOVRSMPLERRCNT          = 16'h0000;    // Offset = 15'h701 Attributes : RO   
parameter L3_RXOVRSMPLERRCNTCLR       = 16'h0000;    // Offset = 15'h702 Attributes : RW   
parameter L3_RXOOBBURST               = 16'h0603;    // Offset = 15'h704 Attributes : RW   
parameter L3_RXOOBCOMINIT             = 16'h2208;    // Offset = 15'h705 Attributes : RW   
parameter L3_RXOOBCOMSAS              = 16'h7525;    // Offset = 15'h706 Attributes : RW   
parameter L3_RXOOBCOMWAKE             = 16'h0603;    // Offset = 15'h707 Attributes : RW   
parameter L3_RXOOBSET                 = 16'h0006;    // Offset = 15'h708 Attributes : RW   
parameter L3_RXOOBSTATUS              = 16'h0000;    // Offset = 15'h709 Attributes : RO   
parameter L3_RXOOBCOMINITCNT          = 16'h0000;    // Offset = 15'h70A Attributes : RO   
parameter L3_RXOOBCOMSASCNT           = 16'h0000;    // Offset = 15'h70B Attributes : RO   
parameter L3_RXOOBCOMWAKECNT          = 16'h0000;    // Offset = 15'h70C Attributes : RO   
parameter L3_RXOOBCNTCLR              = 16'h0000;    // Offset = 15'h70D Attributes : RW   
parameter L3_RXPRBSCHK                = 16'h0001;    // Offset = 15'h710 Attributes : RW   
parameter L3_RXPRBSCHKERRCNT          = 16'h0000;    // Offset = 15'h711 Attributes : RO   
parameter L3_RXPRBSZEROCNT            = 16'h0000;    // Offset = 15'h712 Attributes : RO   
parameter L3_RXPRBSCHKCNTCLR          = 16'h0000;    // Offset = 15'h713 Attributes : RW   
parameter L3_RXPRBSCHKPATTEN1         = 16'h03ff;    // Offset = 15'h714 Attributes : RW   
parameter L3_RXPRBSCHKPATTEN2         = 16'h03ff;    // Offset = 15'h715 Attributes : RW   
parameter L3_RXPRBSCHKPATTEN3         = 16'h0000;    // Offset = 15'h716 Attributes : RW   
parameter L3_RXPRBSCHKPATTEN4         = 16'h0000;    // Offset = 15'h717 Attributes : RW   
parameter L3_RX8B10BCAD               = 16'hc3ff;    // Offset = 15'h720 Attributes : RW   
parameter L3_RX8B10BCADMCOMMA         = 16'h2283;    // Offset = 15'h721 Attributes : RW   
parameter L3_RX8B10BCADPCOMMA         = 16'h217c;    // Offset = 15'h722 Attributes : RW   
parameter L3_RX8B10BCADSLIDE          = 16'h0000;    // Offset = 15'h723 Attributes : RW   
parameter L3_RX8B10BDEC               = 16'h0001;    // Offset = 15'h724 Attributes : RW   
parameter L3_RX8B10BDECCOMMA          = 16'h0000;    // Offset = 15'h725 Attributes : RW   
parameter L3_RX8B10BSYNC              = 16'h5111;    // Offset = 15'h728 Attributes : RW   
parameter L3_RX8B10BSTATUS            = 16'h0000;    // Offset = 15'h729 Attributes : RO   
parameter L3_RX4B5BSET                = 16'h0000;    // Offset = 15'h72B Attributes : RW   
parameter L3_RX4B5BSD                 = 16'h0223;    // Offset = 15'h72C Attributes : RW   
parameter L3_RX4B5BED                 = 16'h0396;    // Offset = 15'h72D Attributes : RW   
parameter L3_RXPMUX                   = 16'h0001;    // Offset = 15'h72F Attributes : RW   
parameter L3_RXLDBUF                  = 16'h0000;    // Offset = 15'h730 Attributes : RW   
parameter L3_RXLDBUFSEQ1              = 16'h0000;    // Offset = 15'h731 Attributes : RW   
parameter L3_RXLDBUFSEQ2              = 16'h0000;    // Offset = 15'h732 Attributes : RW   
parameter L3_RXLDBUFSEQ3              = 16'h0000;    // Offset = 15'h733 Attributes : RW   
parameter L3_RXLDBUFSEQ4              = 16'h0000;    // Offset = 15'h734 Attributes : RW   
parameter L3_RXLDBUFSEQEN             = 16'hf1ff;    // Offset = 15'h735 Attributes : RW   
parameter L3_RXEBUF                   = 16'h0001;    // Offset = 15'h738 Attributes : RW   
parameter L3_RXEBUFCLR                = 16'h0000;    // Offset = 15'h739 Attributes : RW   
parameter L3_RXCLKCOR                 = 16'h0101;    // Offset = 15'h73A Attributes : RW   
parameter L3_RXCLKCORSEQ1             = 16'h011c;    // Offset = 15'h73C Attributes : RW   
parameter L3_RXCLKCORSEQ2             = 16'h0000;    // Offset = 15'h73D Attributes : RW   
parameter L3_RXCLKCORSEQ3             = 16'h0000;    // Offset = 15'h73E Attributes : RW   
parameter L3_RXCLKCORSEQ4             = 16'h0000;    // Offset = 15'h73F Attributes : RW   
parameter L3_RXGEARBOX                = 16'h0000;    // Offset = 15'h740 Attributes : RW   
parameter L3_RXGEARBOXSLIP            = 16'h0000;    // Offset = 15'h741 Attributes : RW   
parameter L3_RXGEARBOXSTATUS          = 16'h0000;    // Offset = 15'h742 Attributes : RO   
parameter L3_RXUIA                    = 16'h0000;    // Offset = 15'h744 Attributes : RW   
parameter L3_PCSCMU                   = 16'hd812;    // Offset = 15'h748 Attributes : RW   
parameter L3_PMAUBRDSET               = 16'h0000;    // Offset = 15'h751 Attributes : RW   
parameter L3_PMAUBRDRSLT              = 16'h0000;    // Offset = 15'h752 Attributes : RO   
parameter L3_PMAUBOFCALSET            = 16'h0000;    // Offset = 15'h753 Attributes : RW   
parameter L3_PMAUBOFCALRSLT           = 16'h0000;    // Offset = 15'h754 Attributes : RO   
parameter L3_PMAUBPHASET              = 16'h0000;    // Offset = 15'h755 Attributes : RW   
parameter L3_PMAUBPHARSLT             = 16'h0000;    // Offset = 15'h756 Attributes : RO   
parameter L3_PCSRMUSRST               = 16'h0000;    // Offset = 15'h758 Attributes : RW   

// PMA CFG Common Regist=ers, Offset = 15'h5000
parameter PMACMU                      = 16'h8e2c;    // Offset = 15'h5000 Attributes : RW   
parameter PMAPLL1                     = 16'h3023;    // Offset = 15'h5001 Attributes : RW   
parameter PMAPLL2                     = 16'h1062;    // Offset = 15'h5002 Attributes : RW   
parameter PMAPLL3                     = 16'h0001;    // Offset = 15'h5003 Attributes : RW   
parameter PMAPLL4                     = 16'h0003;    // Offset = 15'h5004 Attributes : RW   
parameter PMAPLL5                     = 16'h0000;    // Offset = 15'h5005 Attributes : RO   
parameter PMAPLL6                     = 16'h0046;    // Offset = 15'h5006 Attributes : RW   
parameter PMAOSC                      = 16'h00d5;    // Offset = 15'h5007 Attributes : RW   
parameter PMATOP1                     = 16'h8102;    // Offset = 15'h5008 Attributes : RW   
parameter PMATOP2                     = 16'h0002;    // Offset = 15'h5009 Attributes : RW   
parameter PMABG1                      = 16'h0034;    // Offset = 15'h5010 Attributes : RW   
parameter PMABG2                      = 16'h0000;    // Offset = 15'h5011 Attributes : RW   
parameter PMABG3                      = 16'h0000;    // Offset = 15'h5012 Attributes : RW   
parameter PMARESCAL1                  = 16'h0002;    // Offset = 15'h5013 Attributes : RW   
parameter PMARESCAL2                  = 16'h0000;    // Offset = 15'h5014 Attributes : RW   
parameter PMARESCALO1                 = 16'h0000;    // Offset = 15'h5015 Attributes : RO   
parameter PMARESCALO2                 = 16'h0000;    // Offset = 15'h5016 Attributes : RO   
parameter PMARESCAL4                  = 16'h1414;    // Offset = 15'h5017 Attributes : RW   
parameter PMARESCAL5                  = 16'h1414;    // Offset = 15'h5018 Attributes : RW   
parameter PMARESCAL6                  = 16'h0000;    // Offset = 15'h5019 Attributes : RO   
parameter PMAJTAG                     = 16'h000c;    // Offset = 15'h501A Attributes : RW   
parameter PMATOP3                     = 16'h0003;    // Offset = 15'h5020 Attributes : RW   
parameter PMATESTMUX                  = 16'h0000;    // Offset = 15'h5021 Attributes : RW   

// PMA CFG Lane Register=s, Offset = 15'h2000(Lane0) 15'h2200(Lane1) 15'h2400(Lane2) 15'h2600(Lane3) 15'h3000(Broadcast)
parameter L0_TXDRV                    = 16'h400d;    // Offset = 15'h2000 Attributes : RW   
parameter L0_PMATX1                   = 16'h07d4;    // Offset = 15'h2001 Attributes : RW   
parameter L0_PMATX2                   = 16'h3200;    // Offset = 15'h2002 Attributes : RW   
parameter L0_PMATX3                   = 16'h0220;    // Offset = 15'h2003 Attributes : RW   
parameter L0_PMATX4                   = 16'h0008;    // Offset = 15'h2004 Attributes : RW   
parameter L0_PMATX5                   = 16'h0000;    // Offset = 15'h2005 Attributes : RO   
parameter L0_PMATXPHASSC1             = 16'h1d00;    // Offset = 15'h2006 Attributes : RW   
parameter L0_PMATXPHASSC2             = 16'h0000;    // Offset = 15'h2007 Attributes : RW   
parameter L0_PMAACC1                  = 16'h4000;    // Offset = 15'h2008 Attributes : RW   
parameter L0_PMATXPHASSC3             = 16'h0497;    // Offset = 15'h2009 Attributes : RW   
parameter L0_PMARXCDR1                = 16'h2119;    // Offset = 15'h2100 Attributes : RW   
parameter L0_PMARXCDR2                = 16'h071c;    // Offset = 15'h2101 Attributes : RW   
parameter L0_PMARXCDR3                = 16'h2007;    // Offset = 15'h2102 Attributes : RW   
parameter L0_PMARXCDR4                = 16'h1240;    // Offset = 15'h2103 Attributes : RW   
parameter L0_PMARXPHA1                = 16'h0200;    // Offset = 15'h2104 Attributes : RW   
parameter L0_PMARXPHA2                = 16'h0000;    // Offset = 15'h2105 Attributes : RW   
parameter L0_PMARXPHA3                = 16'h0000;    // Offset = 15'h2106 Attributes : RO   
parameter L0_PMARXDEF1                = 16'h9d39;    // Offset = 15'h2107 Attributes : RW   
parameter L0_PMARXDEF2                = 16'h0000;    // Offset = 15'h2108 Attributes : RW   
parameter L0_PMARXDEF3                = 16'h0000;    // Offset = 15'h2109 Attributes : RW   
parameter L0_PMARXDEF4                = 16'h0000;    // Offset = 15'h210A Attributes : RW   
parameter L0_PMARXDEF5                = 16'h0000;    // Offset = 15'h210B Attributes : RO   
parameter L0_PMARXDEF6                = 16'h0000;    // Offset = 15'h210C Attributes : RO   
parameter L0_PMARXDEF7                = 16'h0000;    // Offset = 15'h210D Attributes : RO   
parameter L0_PMARXCTLE1               = 16'h2356;    // Offset = 15'h2110 Attributes : RW   
parameter L0_PMARXCTLE2               = 16'h0000;    // Offset = 15'h2111 Attributes : RO   
parameter L0_PMARXCTLE3               = 16'h0007;    // Offset = 15'h2112 Attributes : RW   
parameter L0_PMARXAFE                 = 16'h005b;    // Offset = 15'h2113 Attributes : RW   
parameter L0_PMARXSQUELCH             = 16'h0031;    // Offset = 15'h2114 Attributes : RW   
parameter L0_PMARXOFCAL1              = 16'h3002;    // Offset = 15'h2115 Attributes : RW   
parameter L0_PMARXOFCAL2              = 16'h0000;    // Offset = 15'h2116 Attributes : RO   
parameter L0_PMARXTOP                 = 16'h0011;    // Offset = 15'h2117 Attributes : RW   

parameter L1_TXDRV                    = 16'h400d;    // Offset = 15'h2200 Attributes : RW   
parameter L1_PMATX1                   = 16'h07d4;    // Offset = 15'h2201 Attributes : RW   
parameter L1_PMATX2                   = 16'h3200;    // Offset = 15'h2202 Attributes : RW   
parameter L1_PMATX3                   = 16'h0220;    // Offset = 15'h2203 Attributes : RW   
parameter L1_PMATX4                   = 16'h0008;    // Offset = 15'h2204 Attributes : RW   
parameter L1_PMATX5                   = 16'h0000;    // Offset = 15'h2205 Attributes : RO   
parameter L1_PMATXPHASSC1             = 16'h1d00;    // Offset = 15'h2206 Attributes : RW   
parameter L1_PMATXPHASSC2             = 16'h0000;    // Offset = 15'h2207 Attributes : RW   
parameter L1_PMAACC1                  = 16'h4000;    // Offset = 15'h2208 Attributes : RW   
parameter L1_PMATXPHASSC3             = 16'h0497;    // Offset = 15'h2209 Attributes : RW   
parameter L1_PMARXCDR1                = 16'h2119;    // Offset = 15'h2300 Attributes : RW   
parameter L1_PMARXCDR2                = 16'h071c;    // Offset = 15'h2301 Attributes : RW   
parameter L1_PMARXCDR3                = 16'h2007;    // Offset = 15'h2302 Attributes : RW   
parameter L1_PMARXCDR4                = 16'h1240;    // Offset = 15'h2303 Attributes : RW   
parameter L1_PMARXPHA1                = 16'h0200;    // Offset = 15'h2304 Attributes : RW   
parameter L1_PMARXPHA2                = 16'h0000;    // Offset = 15'h2305 Attributes : RW   
parameter L1_PMARXPHA3                = 16'h0000;    // Offset = 15'h2306 Attributes : RO   
parameter L1_PMARXDEF1                = 16'h9d39;    // Offset = 15'h2307 Attributes : RW   
parameter L1_PMARXDEF2                = 16'h0000;    // Offset = 15'h2308 Attributes : RW   
parameter L1_PMARXDEF3                = 16'h0000;    // Offset = 15'h2309 Attributes : RW   
parameter L1_PMARXDEF4                = 16'h0000;    // Offset = 15'h230A Attributes : RW   
parameter L1_PMARXDEF5                = 16'h0000;    // Offset = 15'h230B Attributes : RO   
parameter L1_PMARXDEF6                = 16'h0000;    // Offset = 15'h230C Attributes : RO   
parameter L1_PMARXDEF7                = 16'h0000;    // Offset = 15'h230D Attributes : RO   
parameter L1_PMARXCTLE1               = 16'h2356;    // Offset = 15'h2310 Attributes : RW   
parameter L1_PMARXCTLE2               = 16'h0000;    // Offset = 15'h2311 Attributes : RO   
parameter L1_PMARXCTLE3               = 16'h0007;    // Offset = 15'h2312 Attributes : RW   
parameter L1_PMARXAFE                 = 16'h005b;    // Offset = 15'h2313 Attributes : RW   
parameter L1_PMARXSQUELCH             = 16'h0031;    // Offset = 15'h2314 Attributes : RW   
parameter L1_PMARXOFCAL1              = 16'h3002;    // Offset = 15'h2315 Attributes : RW   
parameter L1_PMARXOFCAL2              = 16'h0000;    // Offset = 15'h2316 Attributes : RO   
parameter L1_PMARXTOP                 = 16'h0011;    // Offset = 15'h2317 Attributes : RW   

parameter L2_TXDRV                    = 16'h400d;    // Offset = 15'h2400 Attributes : RW   
parameter L2_PMATX1                   = 16'h07d4;    // Offset = 15'h2401 Attributes : RW   
parameter L2_PMATX2                   = 16'h3200;    // Offset = 15'h2402 Attributes : RW   
parameter L2_PMATX3                   = 16'h0220;    // Offset = 15'h2403 Attributes : RW   
parameter L2_PMATX4                   = 16'h0008;    // Offset = 15'h2404 Attributes : RW   
parameter L2_PMATX5                   = 16'h0000;    // Offset = 15'h2405 Attributes : RO   
parameter L2_PMATXPHASSC1             = 16'h1d00;    // Offset = 15'h2406 Attributes : RW   
parameter L2_PMATXPHASSC2             = 16'h0000;    // Offset = 15'h2407 Attributes : RW   
parameter L2_PMAACC1                  = 16'h4000;    // Offset = 15'h2408 Attributes : RW   
parameter L2_PMATXPHASSC3             = 16'h0497;    // Offset = 15'h2409 Attributes : RW   
parameter L2_PMARXCDR1                = 16'h2119;    // Offset = 15'h2500 Attributes : RW   
parameter L2_PMARXCDR2                = 16'h071c;    // Offset = 15'h2501 Attributes : RW   
parameter L2_PMARXCDR3                = 16'h2007;    // Offset = 15'h2502 Attributes : RW   
parameter L2_PMARXCDR4                = 16'h1240;    // Offset = 15'h2503 Attributes : RW   
parameter L2_PMARXPHA1                = 16'h0200;    // Offset = 15'h2504 Attributes : RW   
parameter L2_PMARXPHA2                = 16'h0000;    // Offset = 15'h2505 Attributes : RW   
parameter L2_PMARXPHA3                = 16'h0000;    // Offset = 15'h2506 Attributes : RO   
parameter L2_PMARXDEF1                = 16'h9d39;    // Offset = 15'h2507 Attributes : RW   
parameter L2_PMARXDEF2                = 16'h0000;    // Offset = 15'h2508 Attributes : RW   
parameter L2_PMARXDEF3                = 16'h0000;    // Offset = 15'h2509 Attributes : RW   
parameter L2_PMARXDEF4                = 16'h0000;    // Offset = 15'h250A Attributes : RW   
parameter L2_PMARXDEF5                = 16'h0000;    // Offset = 15'h250B Attributes : RO   
parameter L2_PMARXDEF6                = 16'h0000;    // Offset = 15'h250C Attributes : RO   
parameter L2_PMARXDEF7                = 16'h0000;    // Offset = 15'h250D Attributes : RO   
parameter L2_PMARXCTLE1               = 16'h2356;    // Offset = 15'h2510 Attributes : RW   
parameter L2_PMARXCTLE2               = 16'h0000;    // Offset = 15'h2511 Attributes : RO   
parameter L2_PMARXCTLE3               = 16'h0007;    // Offset = 15'h2512 Attributes : RW   
parameter L2_PMARXAFE                 = 16'h005b;    // Offset = 15'h2513 Attributes : RW   
parameter L2_PMARXSQUELCH             = 16'h0031;    // Offset = 15'h2514 Attributes : RW   
parameter L2_PMARXOFCAL1              = 16'h3002;    // Offset = 15'h2515 Attributes : RW   
parameter L2_PMARXOFCAL2              = 16'h0000;    // Offset = 15'h2516 Attributes : RO   
parameter L2_PMARXTOP                 = 16'h0011;    // Offset = 15'h2517 Attributes : RW   

parameter L3_TXDRV                    = 16'h400d;    // Offset = 15'h2600 Attributes : RW   
parameter L3_PMATX1                   = 16'h07d4;    // Offset = 15'h2601 Attributes : RW   
parameter L3_PMATX2                   = 16'h3200;    // Offset = 15'h2602 Attributes : RW   
parameter L3_PMATX3                   = 16'h0220;    // Offset = 15'h2603 Attributes : RW   
parameter L3_PMATX4                   = 16'h0008;    // Offset = 15'h2604 Attributes : RW   
parameter L3_PMATX5                   = 16'h0000;    // Offset = 15'h2605 Attributes : RO   
parameter L3_PMATXPHASSC1             = 16'h1d00;    // Offset = 15'h2606 Attributes : RW   
parameter L3_PMATXPHASSC2             = 16'h0000;    // Offset = 15'h2607 Attributes : RW   
parameter L3_PMAACC1                  = 16'h4000;    // Offset = 15'h2608 Attributes : RW   
parameter L3_PMATXPHASSC3             = 16'h0497;    // Offset = 15'h2609 Attributes : RW   
parameter L3_PMARXCDR1                = 16'h2119;    // Offset = 15'h2700 Attributes : RW   
parameter L3_PMARXCDR2                = 16'h071c;    // Offset = 15'h2701 Attributes : RW   
parameter L3_PMARXCDR3                = 16'h2007;    // Offset = 15'h2702 Attributes : RW   
parameter L3_PMARXCDR4                = 16'h1240;    // Offset = 15'h2703 Attributes : RW   
parameter L3_PMARXPHA1                = 16'h0200;    // Offset = 15'h2704 Attributes : RW   
parameter L3_PMARXPHA2                = 16'h0000;    // Offset = 15'h2705 Attributes : RW   
parameter L3_PMARXPHA3                = 16'h0000;    // Offset = 15'h2706 Attributes : RO   
parameter L3_PMARXDEF1                = 16'h9d39;    // Offset = 15'h2707 Attributes : RW   
parameter L3_PMARXDEF2                = 16'h0000;    // Offset = 15'h2708 Attributes : RW   
parameter L3_PMARXDEF3                = 16'h0000;    // Offset = 15'h2709 Attributes : RW   
parameter L3_PMARXDEF4                = 16'h0000;    // Offset = 15'h270A Attributes : RW   
parameter L3_PMARXDEF5                = 16'h0000;    // Offset = 15'h270B Attributes : RO   
parameter L3_PMARXDEF6                = 16'h0000;    // Offset = 15'h270C Attributes : RO   
parameter L3_PMARXDEF7                = 16'h0000;    // Offset = 15'h270D Attributes : RO   
parameter L3_PMARXCTLE1               = 16'h2356;    // Offset = 15'h2710 Attributes : RW   
parameter L3_PMARXCTLE2               = 16'h0000;    // Offset = 15'h2711 Attributes : RO   
parameter L3_PMARXCTLE3               = 16'h0007;    // Offset = 15'h2712 Attributes : RW   
parameter L3_PMARXAFE                 = 16'h005b;    // Offset = 15'h2713 Attributes : RW   
parameter L3_PMARXSQUELCH             = 16'h0031;    // Offset = 15'h2714 Attributes : RW   
parameter L3_PMARXOFCAL1              = 16'h3002;    // Offset = 15'h2715 Attributes : RW   
parameter L3_PMARXOFCAL2              = 16'h0000;    // Offset = 15'h2716 Attributes : RO   
parameter L3_PMARXTOP                 = 16'h0011;    // Offset = 15'h2717 Attributes : RW   

endmodule

module GUC_GPIO (
	rxd_out,
	ted_out,
	txd_out,
	rxd_in,
	ted_in,
	txd_in 
);

output		rxd_out;
output		ted_out;
output		txd_out;
input		rxd_in;
input		ted_in;
input		txd_in;

parameter pd            = 1'b0; 
parameter pu            = 1'b0; 
parameter smt           = 1'b0; 
parameter hv_en         = 1'b0; 
parameter pum           = 8'b0; 
parameter pdm           = 8'b0; 
parameter pdn           = 1'b0; 
parameter odt           = 3'b0; 
parameter gpio_en       = 1'b0; 
parameter jtag_en       = 1'b0; 
parameter drvp          = 3'b0; 
parameter dr3en         = 1'b0; 

mybuf rxd_buf (
	.i	(rxd_in),

	.o	(rxd_out) 
);

mybuf txd_buf (
	.i	(txd_in),

	.o	(txd_out) 
);

mybuf ted_buf (
	.i	(ted_in),

	.o	(ted_out) 
);

endmodule

module mybuf(i,o);

input  i;
output o;

assign o = i;

endmodule
module H6_MAC (
    // Outputs
    a_mac_out, 
    b_mac_out, 
    a_overflow, 
    b_overflow,
    // Inputs
	a_dinxy_cen, b_dinxy_cen,
	a_dinz_cen, b_dinz_cen,
	a_mac_out_cen, b_mac_out_cen,
	a_in_sr, b_in_sr,
	a_out_sr, b_out_sr,
    a_dinx, a_diny, 
    b_dinx, b_diny, 
    a_dinz, b_dinz,
    clk, 
    a_sload, b_sload, 
    a_acc_en, a_dinz_en, 
    b_acc_en, b_dinz_en
);

    //a_mac_out = a_dinx * a_diny + a_dinz;
`ifdef CS_FORMALPRO_HACK
    wire [2:0] modea_sel;
    wire [2:0] modeb_sel;

    wire adinx_input_mode; 
    wire adiny_input_mode; 
    wire adinz_input_mode; 
    wire amac_output_mode; 

    wire bdinx_input_mode; 
    wire bdiny_input_mode; 
    wire bdinz_input_mode; 
    wire bmac_output_mode; 

    wire a_in_rstn_sel;
    wire a_in_setn_sel;
    wire a_sr_syn_sel;
    wire a_ovf_rstn_sel;
    wire [47:0] a_out_rstn_sel;
    wire [47:0] a_out_setn_sel;

    wire b_in_rstn_sel ;
    wire b_in_setn_sel ;
    wire b_sr_syn_sel ;
    wire b_ovf_rstn_sel;
    wire [27:0] b_out_rstn_sel;
    wire [27:0] b_out_setn_sel ;

`else
    parameter modea_sel = 3'b000;
    parameter modeb_sel = 3'b000;

    parameter adinx_input_mode = 1'b0; 
    parameter adiny_input_mode = 1'b0; 
    parameter adinz_input_mode = 1'b0; 
    parameter amac_output_mode = 1'b0; 

    parameter bdinx_input_mode = 1'b0; 
    parameter bdiny_input_mode = 1'b0; 
    parameter bdinz_input_mode = 1'b0; 
    parameter bmac_output_mode = 1'b0; 

    parameter a_in_rstn_sel = 1'b0;
    parameter a_in_setn_sel = 1'b0;
    parameter a_sr_syn_sel= 1'b0;
    parameter a_ovf_rstn_sel= 1'b0;
    parameter [47:0] a_out_rstn_sel= 48'b0;
    parameter [47:0] a_out_setn_sel= 48'b0;
    parameter a_out_rstn_sel_h = 24'b0;
    parameter a_out_rstn_sel_l = 24'b0;
    parameter a_out_setn_sel_h = 24'b0;
    parameter a_out_setn_sel_l = 24'b0;

    parameter b_in_rstn_sel = 1'b0;
    parameter b_in_setn_sel = 1'b0;
    parameter b_sr_syn_sel= 1'b0;
    parameter b_ovf_rstn_sel= 1'b0;
    parameter b_out_rstn_sel= 28'b0;
    parameter b_out_setn_sel= 28'b0;
`endif

//---------------------------------------------------------------------------------
//for SW
//---------------------------------------------------------------------------------
    //parameter modea_sel = ""; //"18x18", "12x9", "9x9"
    //parameter modeb_sel = ""; //"18x18", "12x9", "9x9"

    //parameter adinx_input_mode = "bypass"; //"register" 
    //parameter adiny_input_mode = "bypass"; //"register" 
    //parameter adinz_input_mode = "bypass"; //"register" 
    //parameter amac_output_mode = "bypass"; //"register" 

    //parameter bdinx_input_mode = "bypass"; //"register" 
    //parameter bdiny_input_mode = "bypass"; //"register" 
    //parameter bdinz_input_mode = "bypass"; //"register" 
    //parameter bmac_output_mode = "bypass"; //"register" 
//---------------------------------------------------------------------------------

	input	a_dinxy_cen, b_dinxy_cen;
	input	a_dinz_cen, b_dinz_cen;
	input	a_mac_out_cen, b_mac_out_cen;
	input	a_in_sr, b_in_sr;
	input	a_out_sr, b_out_sr;

    //Group A, multiplier input
    input [13:0] a_dinx ;
    input [9:0]  a_diny ;
    
    //Group B, multiplier input
    input [13:0] b_dinx ;
    input [9:0]  b_diny ;
    
    //Group A,B, post add input
    input [24:0] a_dinz;
    input [24:0] b_dinz;
    
    //global signal
    input clk;
    
    //acculate load 
    input a_sload;
    input b_sload;
    
    //acculate en
    input a_acc_en;
    input b_acc_en;
    
    //post add en
    input a_dinz_en;
    input b_dinz_en;
    
    //Group A,B multiplier/acculate output
    output [24:0] a_mac_out;
    output [24:0] b_mac_out;
    
    //Group A,B overflow
    output a_overflow;
    output b_overflow;

	wire clk_in;
	wire rstn_in;
	
	//a mac
	wire [12:0] a_x_in ;
	wire [9:0]  a_y_in ;
	wire [24:0] a_z_in;
	
	reg [12:0] a_qx_o_mux ;
	reg [12:0] a_qx_o_reg_syn ;
	reg [12:0] a_qx_o_reg_asyn ;
	wire [12:0] a_qx_o_reg ;
	
	reg [9:0] a_qy_o_mux ;
	reg [9:0] a_qy_o_reg_syn ;
	reg [9:0] a_qy_o_reg_asyn ;
	wire [9:0] a_qy_o_reg ;
	
	reg [24:0] a_qz_o_mux ;
	reg [24:0] a_qz_o_reg_syn ;
	reg [24:0] a_qz_o_reg_asyn ;
	wire [24:0] a_qz_o_reg ;
	
	wire [24:0] a_mult_o ;
	wire [24:0] a_qmac_o_reg;
	wire [24:0] a_qmac_i;
	wire  [24:0] a_qmac_o_reg_syn;
	wire  [24:0] a_qmac_o_reg_asyn;
	reg [24:0] a_add_mux ;
	wire [24:0] a_mac_o_mux ;
	wire [24:0] a_mac_o_out ;
	wire [24:0] a_add_o ;

	wire mac_a_overflow;
	wire a_overflow_tmp;
	wire b_overflow_tmp;
	wire mac_overflow_tmp;//for 18x18
	wire mac_overflow;//for 18x18

    wire  mac_a_overflow_d;
    reg   mac_a_overflow_d_asyn;
    reg   mac_a_overflow_d_syn;
	reg   mac_a_overflow_temp_asyn ;
	wire  mac_a_overflow_or ;
    wire  mac_b_overflow_d;
    reg   mac_b_overflow_d_asyn;
    reg   mac_b_overflow_d_syn;
	reg   mac_b_overflow_temp_asyn ;
	wire  mac_b_overflow_or ;
	reg   mac_overflow_d_asyn;//for 18x18
	reg   mac_overflow_d_syn;//for 18x18
	reg   mac_overflow_temp_asyn ;//for 18x18
	wire  mac_overflow_or ;//for 18x18
	wire  mac_overflow_d;//for 18x18
		
	wire a_signedx;
	wire a_signedy;
	wire a_signedz;
	
	wire a_sload_i;
	wire a_acc_en_i; 
    reg  a_dinz_en_i;
    wire  a_dinz_en_reg;
    reg  a_dinz_en_reg_asyn;
    reg  a_dinz_en_reg_syn;

	wire a_in_rstn ;
	wire a_in_setn ;
	wire a_ovf_rstn;
	wire a_0_out_rstn;
	wire a_1_out_rstn;
	wire a_2_out_rstn;
	wire a_3_out_rstn;
	wire a_4_out_rstn;
	wire a_5_out_rstn;
	wire a_6_out_rstn;
	wire a_7_out_rstn;
	wire a_8_out_rstn;
	wire a_9_out_rstn;
	wire a_10_out_rstn;
	wire a_11_out_rstn;
	wire a_12_out_rstn;
	wire a_13_out_rstn;
	wire a_14_out_rstn;
	wire a_15_out_rstn;
	wire a_16_out_rstn;
	wire a_17_out_rstn;
	wire a_18_out_rstn;
	wire a_19_out_rstn;
	wire a_20_out_rstn;
	wire a_21_out_rstn;
	wire a_22_out_rstn;
	wire a_23_out_rstn;
	wire a_24_out_rstn;
	wire a_25_out_rstn;
	wire a_26_out_rstn;
	wire a_27_out_rstn;
	wire a_28_out_rstn;
	wire a_29_out_rstn;
	wire a_30_out_rstn;
	wire a_31_out_rstn;
	wire a_32_out_rstn;
	wire a_33_out_rstn;
	wire a_34_out_rstn;
	wire a_35_out_rstn;
	wire a_36_out_rstn;
	wire a_37_out_rstn;
	wire a_38_out_rstn;
	wire a_39_out_rstn;
	wire a_40_out_rstn;
	wire a_41_out_rstn;
	wire a_42_out_rstn;
	wire a_43_out_rstn;
	wire a_44_out_rstn;
	wire a_45_out_rstn;
	wire a_46_out_rstn;
	wire a_47_out_rstn;

	wire a_0_out_setn;
	wire a_1_out_setn;
	wire a_2_out_setn;
	wire a_3_out_setn;
	wire a_4_out_setn;
	wire a_5_out_setn;
	wire a_6_out_setn;
	wire a_7_out_setn;
	wire a_8_out_setn;
	wire a_9_out_setn;
	wire a_10_out_setn;
	wire a_11_out_setn;
	wire a_12_out_setn;
	wire a_13_out_setn;
	wire a_14_out_setn;
	wire a_15_out_setn;
	wire a_16_out_setn;
	wire a_17_out_setn;
	wire a_18_out_setn;
	wire a_19_out_setn;
	wire a_20_out_setn;
	wire a_21_out_setn;
	wire a_22_out_setn;
	wire a_23_out_setn;
	wire a_24_out_setn;
	wire a_25_out_setn;
	wire a_26_out_setn;
	wire a_27_out_setn;
	wire a_28_out_setn;
	wire a_29_out_setn;
	wire a_30_out_setn;
	wire a_31_out_setn;
	wire a_32_out_setn;
	wire a_33_out_setn;
	wire a_34_out_setn;
	wire a_35_out_setn;
	wire a_36_out_setn;
	wire a_37_out_setn;
	wire a_38_out_setn;
	wire a_39_out_setn;
	wire a_40_out_setn;
	wire a_41_out_setn;
	wire a_42_out_setn;
	wire a_43_out_setn;
	wire a_44_out_setn;
	wire a_45_out_setn;
	wire a_46_out_setn;
	wire a_47_out_setn;
	
	wire b_in_rstn ;
	wire b_in_setn ;
	wire b_ovf_rstn ;
	wire b_0_out_rstn;
	wire b_1_out_rstn;
	wire b_2_out_rstn;
	wire b_3_out_rstn;
	wire b_4_out_rstn;
	wire b_5_out_rstn;
	wire b_6_out_rstn;
	wire b_7_out_rstn;
	wire b_8_out_rstn;
	wire b_9_out_rstn;
	wire b_10_out_rstn;
	wire b_11_out_rstn;
	wire b_12_out_rstn;
	wire b_13_out_rstn;
	wire b_14_out_rstn;
	wire b_15_out_rstn;
	wire b_16_out_rstn;
	wire b_17_out_rstn;
	wire b_18_out_rstn;
	wire b_19_out_rstn;
	wire b_20_out_rstn;
	wire b_21_out_rstn;
	wire b_22_out_rstn;
	wire b_23_out_rstn;
	wire b_24_out_rstn;

	wire b_0_out_setn;
	wire b_1_out_setn;
	wire b_2_out_setn;
	wire b_3_out_setn;
	wire b_4_out_setn;
	wire b_5_out_setn;
	wire b_6_out_setn;
	wire b_7_out_setn;
	wire b_8_out_setn;
	wire b_9_out_setn;
	wire b_10_out_setn;
	wire b_11_out_setn;
	wire b_12_out_setn;
	wire b_13_out_setn;
	wire b_14_out_setn;
	wire b_15_out_setn;
	wire b_16_out_setn;
	wire b_17_out_setn;
	wire b_18_out_setn;
	wire b_19_out_setn;
	wire b_20_out_setn;
	wire b_21_out_setn;
	wire b_22_out_setn;
	wire b_23_out_setn;
	wire b_24_out_setn;
//generate set/reset signal
assign a_in_rstn  = a_in_rstn_sel  == 1 ? a_in_sr : 1'b1;
assign a_in_setn  = a_in_setn_sel  == 1 ? a_in_sr : 1'b1;
assign a_ovf_rstn = a_ovf_rstn_sel == 1 ? a_out_sr : 1'b1;
assign a_0_out_rstn = a_out_rstn_sel[0] == 1 ? a_out_sr : 1'b1;
assign a_1_out_rstn = a_out_rstn_sel[1] == 1 ? a_out_sr : 1'b1;
assign a_2_out_rstn = a_out_rstn_sel[2] == 1 ? a_out_sr : 1'b1;
assign a_3_out_rstn = a_out_rstn_sel[3] == 1 ? a_out_sr : 1'b1;
assign a_4_out_rstn = a_out_rstn_sel[4] == 1 ? a_out_sr : 1'b1;
assign a_5_out_rstn = a_out_rstn_sel[5] == 1 ? a_out_sr : 1'b1;
assign a_6_out_rstn = a_out_rstn_sel[6] == 1 ? a_out_sr : 1'b1;
assign a_7_out_rstn = a_out_rstn_sel[7] == 1 ? a_out_sr : 1'b1;
assign a_8_out_rstn = a_out_rstn_sel[8] == 1 ? a_out_sr : 1'b1;
assign a_9_out_rstn = a_out_rstn_sel[9] == 1 ? a_out_sr : 1'b1;
assign a_10_out_rstn = a_out_rstn_sel[10] == 1 ? a_out_sr : 1'b1;
assign a_11_out_rstn = a_out_rstn_sel[11] == 1 ? a_out_sr : 1'b1;
assign a_12_out_rstn = a_out_rstn_sel[12] == 1 ? a_out_sr : 1'b1;
assign a_13_out_rstn = a_out_rstn_sel[13] == 1 ? a_out_sr : 1'b1;
assign a_14_out_rstn = a_out_rstn_sel[14] == 1 ? a_out_sr : 1'b1;
assign a_15_out_rstn = a_out_rstn_sel[15] == 1 ? a_out_sr : 1'b1;
assign a_16_out_rstn = a_out_rstn_sel[16] == 1 ? a_out_sr : 1'b1;
assign a_17_out_rstn = a_out_rstn_sel[17] == 1 ? a_out_sr : 1'b1;
assign a_18_out_rstn = a_out_rstn_sel[18] == 1 ? a_out_sr : 1'b1;
assign a_19_out_rstn = a_out_rstn_sel[19] == 1 ? a_out_sr : 1'b1;
assign a_20_out_rstn = a_out_rstn_sel[20] == 1 ? a_out_sr : 1'b1;
assign a_21_out_rstn = a_out_rstn_sel[21] == 1 ? a_out_sr : 1'b1;
assign a_22_out_rstn = a_out_rstn_sel[22] == 1 ? a_out_sr : 1'b1;
assign a_23_out_rstn = a_out_rstn_sel[23] == 1 ? a_out_sr : 1'b1;
assign a_24_out_rstn = a_out_rstn_sel[24] == 1 ? a_out_sr : 1'b1;
assign a_25_out_rstn = a_out_rstn_sel[25] == 1 ? a_out_sr : 1'b1;
assign a_26_out_rstn = a_out_rstn_sel[26] == 1 ? a_out_sr : 1'b1;
assign a_27_out_rstn = a_out_rstn_sel[27] == 1 ? a_out_sr : 1'b1;
assign a_28_out_rstn = a_out_rstn_sel[28] == 1 ? a_out_sr : 1'b1;
assign a_29_out_rstn = a_out_rstn_sel[29] == 1 ? a_out_sr : 1'b1;
assign a_30_out_rstn = a_out_rstn_sel[30] == 1 ? a_out_sr : 1'b1;
assign a_31_out_rstn = a_out_rstn_sel[31] == 1 ? a_out_sr : 1'b1;
assign a_32_out_rstn = a_out_rstn_sel[32] == 1 ? a_out_sr : 1'b1;
assign a_33_out_rstn = a_out_rstn_sel[33] == 1 ? a_out_sr : 1'b1;
assign a_34_out_rstn = a_out_rstn_sel[34] == 1 ? a_out_sr : 1'b1;
assign a_35_out_rstn = a_out_rstn_sel[35] == 1 ? a_out_sr : 1'b1;
assign a_36_out_rstn = a_out_rstn_sel[36] == 1 ? a_out_sr : 1'b1;
assign a_37_out_rstn = a_out_rstn_sel[37] == 1 ? a_out_sr : 1'b1;
assign a_38_out_rstn = a_out_rstn_sel[38] == 1 ? a_out_sr : 1'b1;
assign a_39_out_rstn = a_out_rstn_sel[39] == 1 ? a_out_sr : 1'b1;
assign a_40_out_rstn = a_out_rstn_sel[40] == 1 ? a_out_sr : 1'b1;
assign a_41_out_rstn = a_out_rstn_sel[41] == 1 ? a_out_sr : 1'b1;
assign a_42_out_rstn = a_out_rstn_sel[42] == 1 ? a_out_sr : 1'b1;
assign a_43_out_rstn = a_out_rstn_sel[43] == 1 ? a_out_sr : 1'b1;
assign a_44_out_rstn = a_out_rstn_sel[44] == 1 ? a_out_sr : 1'b1;
assign a_45_out_rstn = a_out_rstn_sel[45] == 1 ? a_out_sr : 1'b1;
assign a_46_out_rstn = a_out_rstn_sel[46] == 1 ? a_out_sr : 1'b1;
assign a_47_out_rstn = a_out_rstn_sel[47] == 1 ? a_out_sr : 1'b1;

assign a_0_out_setn = a_out_setn_sel[0] == 1 ? a_out_sr : 1'b1;
assign a_1_out_setn = a_out_setn_sel[1] == 1 ? a_out_sr : 1'b1;
assign a_2_out_setn = a_out_setn_sel[2] == 1 ? a_out_sr : 1'b1;
assign a_3_out_setn = a_out_setn_sel[3] == 1 ? a_out_sr : 1'b1;
assign a_4_out_setn = a_out_setn_sel[4] == 1 ? a_out_sr : 1'b1;
assign a_5_out_setn = a_out_setn_sel[5] == 1 ? a_out_sr : 1'b1;
assign a_6_out_setn = a_out_setn_sel[6] == 1 ? a_out_sr : 1'b1;
assign a_7_out_setn = a_out_setn_sel[7] == 1 ? a_out_sr : 1'b1;
assign a_8_out_setn = a_out_setn_sel[8] == 1 ? a_out_sr : 1'b1;
assign a_9_out_setn = a_out_setn_sel[9] == 1 ? a_out_sr : 1'b1;
assign a_10_out_setn = a_out_setn_sel[10] == 1 ? a_out_sr : 1'b1;
assign a_11_out_setn = a_out_setn_sel[11] == 1 ? a_out_sr : 1'b1;
assign a_12_out_setn = a_out_setn_sel[12] == 1 ? a_out_sr : 1'b1;
assign a_13_out_setn = a_out_setn_sel[13] == 1 ? a_out_sr : 1'b1;
assign a_14_out_setn = a_out_setn_sel[14] == 1 ? a_out_sr : 1'b1;
assign a_15_out_setn = a_out_setn_sel[15] == 1 ? a_out_sr : 1'b1;
assign a_16_out_setn = a_out_setn_sel[16] == 1 ? a_out_sr : 1'b1;
assign a_17_out_setn = a_out_setn_sel[17] == 1 ? a_out_sr : 1'b1;
assign a_18_out_setn = a_out_setn_sel[18] == 1 ? a_out_sr : 1'b1;
assign a_19_out_setn = a_out_setn_sel[19] == 1 ? a_out_sr : 1'b1;
assign a_20_out_setn = a_out_setn_sel[20] == 1 ? a_out_sr : 1'b1;
assign a_21_out_setn = a_out_setn_sel[21] == 1 ? a_out_sr : 1'b1;
assign a_22_out_setn = a_out_setn_sel[22] == 1 ? a_out_sr : 1'b1;
assign a_23_out_setn = a_out_setn_sel[23] == 1 ? a_out_sr : 1'b1;
assign a_24_out_setn = a_out_setn_sel[24] == 1 ? a_out_sr : 1'b1;
assign a_25_out_setn = a_out_setn_sel[25] == 1 ? a_out_sr : 1'b1;
assign a_26_out_setn = a_out_setn_sel[26] == 1 ? a_out_sr : 1'b1;
assign a_27_out_setn = a_out_setn_sel[27] == 1 ? a_out_sr : 1'b1;
assign a_28_out_setn = a_out_setn_sel[28] == 1 ? a_out_sr : 1'b1;
assign a_29_out_setn = a_out_setn_sel[29] == 1 ? a_out_sr : 1'b1;
assign a_30_out_setn = a_out_setn_sel[30] == 1 ? a_out_sr : 1'b1;
assign a_31_out_setn = a_out_setn_sel[31] == 1 ? a_out_sr : 1'b1;
assign a_32_out_setn = a_out_setn_sel[32] == 1 ? a_out_sr : 1'b1;
assign a_33_out_setn = a_out_setn_sel[33] == 1 ? a_out_sr : 1'b1;
assign a_34_out_setn = a_out_setn_sel[34] == 1 ? a_out_sr : 1'b1;
assign a_35_out_setn = a_out_setn_sel[35] == 1 ? a_out_sr : 1'b1;
assign a_36_out_setn = a_out_setn_sel[36] == 1 ? a_out_sr : 1'b1;
assign a_37_out_setn = a_out_setn_sel[37] == 1 ? a_out_sr : 1'b1;
assign a_38_out_setn = a_out_setn_sel[38] == 1 ? a_out_sr : 1'b1;
assign a_39_out_setn = a_out_setn_sel[39] == 1 ? a_out_sr : 1'b1;
assign a_40_out_setn = a_out_setn_sel[40] == 1 ? a_out_sr : 1'b1;
assign a_41_out_setn = a_out_setn_sel[41] == 1 ? a_out_sr : 1'b1;
assign a_42_out_setn = a_out_setn_sel[42] == 1 ? a_out_sr : 1'b1;
assign a_43_out_setn = a_out_setn_sel[43] == 1 ? a_out_sr : 1'b1;
assign a_44_out_setn = a_out_setn_sel[44] == 1 ? a_out_sr : 1'b1;
assign a_45_out_setn = a_out_setn_sel[45] == 1 ? a_out_sr : 1'b1;
assign a_46_out_setn = a_out_setn_sel[46] == 1 ? a_out_sr : 1'b1;
assign a_47_out_setn = a_out_setn_sel[47] == 1 ? a_out_sr : 1'b1;

assign b_in_rstn  = b_in_rstn_sel  == 1 ? b_in_sr : 1'b1;
assign b_in_setn  = b_in_setn_sel  == 1 ? b_in_sr : 1'b1;
assign b_ovf_rstn = b_ovf_rstn_sel == 1 ? b_out_sr : 1'b1;
assign b_0_out_rstn = b_out_rstn_sel[0] == 1 ? b_out_sr : 1'b1;
assign b_1_out_rstn = b_out_rstn_sel[1] == 1 ? b_out_sr : 1'b1;
assign b_2_out_rstn = b_out_rstn_sel[2] == 1 ? b_out_sr : 1'b1;
assign b_3_out_rstn = b_out_rstn_sel[3] == 1 ? b_out_sr : 1'b1;
assign b_4_out_rstn = b_out_rstn_sel[4] == 1 ? b_out_sr : 1'b1;
assign b_5_out_rstn = b_out_rstn_sel[5] == 1 ? b_out_sr : 1'b1;
assign b_6_out_rstn = b_out_rstn_sel[6] == 1 ? b_out_sr : 1'b1;
assign b_7_out_rstn = b_out_rstn_sel[7] == 1 ? b_out_sr : 1'b1;
assign b_8_out_rstn = b_out_rstn_sel[8] == 1 ? b_out_sr : 1'b1;
assign b_9_out_rstn = b_out_rstn_sel[9] == 1 ? b_out_sr : 1'b1;
assign b_10_out_rstn = b_out_rstn_sel[10] == 1 ? b_out_sr : 1'b1;
assign b_11_out_rstn = b_out_rstn_sel[11] == 1 ? b_out_sr : 1'b1;
assign b_12_out_rstn = b_out_rstn_sel[12] == 1 ? b_out_sr : 1'b1;
assign b_13_out_rstn = b_out_rstn_sel[13] == 1 ? b_out_sr : 1'b1;
assign b_14_out_rstn = b_out_rstn_sel[14] == 1 ? b_out_sr : 1'b1;
assign b_15_out_rstn = b_out_rstn_sel[15] == 1 ? b_out_sr : 1'b1;
assign b_16_out_rstn = b_out_rstn_sel[16] == 1 ? b_out_sr : 1'b1;
assign b_17_out_rstn = b_out_rstn_sel[17] == 1 ? b_out_sr : 1'b1;
assign b_18_out_rstn = b_out_rstn_sel[18] == 1 ? b_out_sr : 1'b1;
assign b_19_out_rstn = b_out_rstn_sel[19] == 1 ? b_out_sr : 1'b1;
assign b_20_out_rstn = b_out_rstn_sel[20] == 1 ? b_out_sr : 1'b1;
assign b_21_out_rstn = b_out_rstn_sel[21] == 1 ? b_out_sr : 1'b1;
assign b_22_out_rstn = b_out_rstn_sel[22] == 1 ? b_out_sr : 1'b1;
assign b_23_out_rstn = b_out_rstn_sel[23] == 1 ? b_out_sr : 1'b1;
assign b_24_out_rstn = b_out_rstn_sel[24] == 1 ? b_out_sr : 1'b1;

assign b_0_out_setn = b_out_setn_sel[0] == 1 ? b_out_sr : 1'b1;
assign b_1_out_setn = b_out_setn_sel[1] == 1 ? b_out_sr : 1'b1;
assign b_2_out_setn = b_out_setn_sel[2] == 1 ? b_out_sr : 1'b1;
assign b_3_out_setn = b_out_setn_sel[3] == 1 ? b_out_sr : 1'b1;
assign b_4_out_setn = b_out_setn_sel[4] == 1 ? b_out_sr : 1'b1;
assign b_5_out_setn = b_out_setn_sel[5] == 1 ? b_out_sr : 1'b1;
assign b_6_out_setn = b_out_setn_sel[6] == 1 ? b_out_sr : 1'b1;
assign b_7_out_setn = b_out_setn_sel[7] == 1 ? b_out_sr : 1'b1;
assign b_8_out_setn = b_out_setn_sel[8] == 1 ? b_out_sr : 1'b1;
assign b_9_out_setn = b_out_setn_sel[9] == 1 ? b_out_sr : 1'b1;
assign b_10_out_setn = b_out_setn_sel[10] == 1 ? b_out_sr : 1'b1;
assign b_11_out_setn = b_out_setn_sel[11] == 1 ? b_out_sr : 1'b1;
assign b_12_out_setn = b_out_setn_sel[12] == 1 ? b_out_sr : 1'b1;
assign b_13_out_setn = b_out_setn_sel[13] == 1 ? b_out_sr : 1'b1;
assign b_14_out_setn = b_out_setn_sel[14] == 1 ? b_out_sr : 1'b1;
assign b_15_out_setn = b_out_setn_sel[15] == 1 ? b_out_sr : 1'b1;
assign b_16_out_setn = b_out_setn_sel[16] == 1 ? b_out_sr : 1'b1;
assign b_17_out_setn = b_out_setn_sel[17] == 1 ? b_out_sr : 1'b1;
assign b_18_out_setn = b_out_setn_sel[18] == 1 ? b_out_sr : 1'b1;
assign b_19_out_setn = b_out_setn_sel[19] == 1 ? b_out_sr : 1'b1;
assign b_20_out_setn = b_out_setn_sel[20] == 1 ? b_out_sr : 1'b1;
assign b_21_out_setn = b_out_setn_sel[21] == 1 ? b_out_sr : 1'b1;
assign b_22_out_setn = b_out_setn_sel[22] == 1 ? b_out_sr : 1'b1;
assign b_23_out_setn = b_out_setn_sel[23] == 1 ? b_out_sr : 1'b1;
assign b_24_out_setn = b_out_setn_sel[24] == 1 ? b_out_sr : 1'b1;
	
	wire a_xreg = (adinx_input_mode == "register") || (adinx_input_mode == 1); 
	wire a_yreg = (adiny_input_mode == "register") || (adiny_input_mode == 1); 
	wire a_zreg = (adinz_input_mode == "register") || (adinz_input_mode == 1); 
	wire a_macreg = (amac_output_mode == "register") || (amac_output_mode == 1); 	
		
	//b mac
	wire [12:0] b_x_in ;
	wire [9:0]  b_y_in ;
	wire [24:0] b_z_in;
	
	reg [12:0] b_qx_o_mux ;
	wire [12:0] b_qx_o_reg ;
	reg  [12:0] b_qx_o_reg_asyn ;
	reg  [12:0] b_qx_o_reg_syn ;
	
	reg [9:0] b_qy_o_mux ;
	wire [9:0] b_qy_o_reg ;
	reg [9:0] b_qy_o_reg_asyn ;
	reg [9:0] b_qy_o_reg_syn ;
	
	reg [24:0] b_qz_o_mux ;
	wire [24:0] b_qz_o_reg ;
	reg [24:0] b_qz_o_reg_asyn ;
	reg [24:0] b_qz_o_reg_syn ;
	
	wire [24:0] b_mult_o ;
	wire [24:0] b_qmac_o_reg_asyn;
	wire [24:0] b_qmac_o_reg_syn;
	wire [24:0] b_qmac_o_reg;
	wire [24:0] b_qmac_i ;
	reg [24:0] b_add_mux ;
	wire [24:0] b_mac_o_mux ;
	wire [24:0] b_mac_o_out ;
	wire [24:0] b_add_o ;
		
	wire b_signedx;
	wire b_signedy;
	wire b_signedz;
	
	wire b_sload_i;
	wire b_acc_en_i; 
    reg  b_dinz_en_i;
    wire  b_dinz_en_reg;
    reg  b_dinz_en_reg_asyn;
    reg  b_dinz_en_reg_syn;
	
	wire b_xreg = (bdinx_input_mode == "register") || (bdinx_input_mode == 1); 
	wire b_yreg = (bdiny_input_mode == "register") || (bdiny_input_mode == 1); 
	wire b_zreg = (bdinz_input_mode == "register") || (bdinz_input_mode == 1); 
	wire b_macreg = (bmac_output_mode == "register") || (bmac_output_mode == 1); 
		
	//18x18 mac
	wire [17:0] x_in ;
	wire [17:0] y_in ;
	wire [47:0] z_in;
	
	wire [17:0] qx_o_mux ;
	
	wire [17:0] qy_o_mux ;
	
	wire [47:0] qz_o_mux ;
	
	wire [47:0] mult_o ;
	wire [47:0]  qmac_o_reg_asyn;
	wire [47:0]  qmac_o_reg_syn;
	wire [47:0] qmac_o_reg;
	wire [47:0] qmac_i;
	reg [47:0] add_mux ;
	wire [47:0] mac_o_mux ;
	wire [47:0] add_o ;
		
	wire signedx;
	wire signedy;
	wire signedz;
	
	wire sload_i;
	wire acc_en_i, dinz_en_i;
	
	wire xreg =   (adinx_input_mode == "register") || (adinx_input_mode == 1); 
	wire yreg =   (adiny_input_mode == "register") || (adiny_input_mode == 1); 
	wire zreg =   (adinz_input_mode == "register") || (adinz_input_mode == 1); 
	wire macreg = (amac_output_mode == "register") || (amac_output_mode == 1); 
	
	assign signedx = b_signedx;
	assign signedy = b_signedy;
	//assign signedz = b_z_in[19 ];
	assign signedz = b_qz_o_mux[23];
	
	assign sload_i = a_sload_i;
	assign acc_en_i = a_acc_en_i;
	assign dinz_en_i = a_dinz_en_i;
	
	buf b_clk (clk_in, clk);
		  
	//buf b_a_signedx	(a_signedx, a_dinx[13]);
	//buf b_a_signedy	(a_signedy, a_diny[9]);
	//buf b_a_signedz	(a_signedz, a_dinz[20]);
    assign a_signedx = a_qx_o_mux[12];
    assign a_signedy = a_qy_o_mux[9];
    assign a_signedz = a_qz_o_mux[24];
	   
	buf b_a_x_in_0 	(a_x_in[0 ], a_dinx[0 ]);
	buf b_a_x_in_1 	(a_x_in[1 ], a_dinx[1 ]);
	buf b_a_x_in_2 	(a_x_in[2 ], a_dinx[2 ]);
	buf b_a_x_in_3 	(a_x_in[3 ], a_dinx[3 ]);
	buf b_a_x_in_4 	(a_x_in[4 ], a_dinx[4 ]);
	buf b_a_x_in_5 	(a_x_in[5 ], a_dinx[5 ]);
	buf b_a_x_in_6 	(a_x_in[6 ], a_dinx[6 ]);
	buf b_a_x_in_7 	(a_x_in[7 ], a_dinx[7 ]);
	buf b_a_x_in_8 	(a_x_in[8 ], a_dinx[8 ]);
	buf b_a_x_in_9 	(a_x_in[9 ], a_dinx[9 ]);
	buf b_a_x_in_10 (a_x_in[10], a_dinx[10]);
	buf b_a_x_in_11 (a_x_in[11], a_dinx[11]);	
	buf b_a_x_in_12 (a_x_in[12], a_dinx[12]);	
	    
	buf b_a_y_in_0 	(a_y_in[0 ], a_diny[0 ]);
	buf b_a_y_in_1 	(a_y_in[1 ], a_diny[1 ]);
	buf b_a_y_in_2 	(a_y_in[2 ], a_diny[2 ]);
	buf b_a_y_in_3 	(a_y_in[3 ], a_diny[3 ]);
	buf b_a_y_in_4 	(a_y_in[4 ], a_diny[4 ]);
	buf b_a_y_in_5 	(a_y_in[5 ], a_diny[5 ]);
	buf b_a_y_in_6 	(a_y_in[6 ], a_diny[6 ]);
	buf b_a_y_in_7 	(a_y_in[7 ], a_diny[7 ]);
	buf b_a_y_in_8 	(a_y_in[8 ], a_diny[8 ]);
	buf b_a_y_in_9 	(a_y_in[9 ], a_diny[9 ]);
	   
	buf b_a_z_in_0 	(a_z_in[0  ], a_dinz[0 ]);
	buf b_a_z_in_1 	(a_z_in[1  ], a_dinz[1 ]);
	buf b_a_z_in_2 	(a_z_in[2  ], a_dinz[2 ]);
	buf b_a_z_in_3 	(a_z_in[3  ], a_dinz[3 ]);
	buf b_a_z_in_4 	(a_z_in[4  ], a_dinz[4 ]);
	buf b_a_z_in_5 	(a_z_in[5  ], a_dinz[5 ]);
	buf b_a_z_in_6 	(a_z_in[6  ], a_dinz[6 ]);
	buf b_a_z_in_7 	(a_z_in[7  ], a_dinz[7 ]);
	buf b_a_z_in_8 	(a_z_in[8  ], a_dinz[8 ]);
	buf b_a_z_in_9 	(a_z_in[9  ], a_dinz[9 ]);
	buf b_a_z_in_10 (a_z_in[10 ], a_dinz[10]);
	buf b_a_z_in_11 (a_z_in[11 ], a_dinz[11]);	
	buf b_a_z_in_12 (a_z_in[12 ], a_dinz[12]);
	buf b_a_z_in_13 (a_z_in[13 ], a_dinz[13]);
	buf b_a_z_in_14 (a_z_in[14 ], a_dinz[14]);
	buf b_a_z_in_15 (a_z_in[15 ], a_dinz[15]);
	buf b_a_z_in_16 (a_z_in[16 ], a_dinz[16]);
	buf b_a_z_in_17 (a_z_in[17 ], a_dinz[17]);
	buf b_a_z_in_18 (a_z_in[18 ], a_dinz[18]);
	buf b_a_z_in_19 (a_z_in[19 ], a_dinz[19]);
	buf b_a_z_in_20 (a_z_in[20 ], a_dinz[20]);
	buf b_a_z_in_21 (a_z_in[21 ], a_dinz[21]);
	buf b_a_z_in_22 (a_z_in[22 ], a_dinz[22]);
	buf b_a_z_in_23 (a_z_in[23 ], a_dinz[23]);
	buf b_a_z_in_24 (a_z_in[24 ], a_dinz[24]);
	
	//buf b_b_signedx (b_signedx, b_dinx[13]);
	//buf b_b_signedy (b_signedy, b_diny[9]);
	//buf b_b_signedz (b_signedz, b_dinz[20]);
    assign b_signedx = b_qx_o_mux[12];
    assign b_signedy = b_qy_o_mux[9];
    assign b_signedz = b_qz_o_mux[24];
	    
	buf b_b_x_in_0 	(b_x_in[0 ], b_dinx[0 ]);
	buf b_b_x_in_1 	(b_x_in[1 ], b_dinx[1 ]);
	buf b_b_x_in_2 	(b_x_in[2 ], b_dinx[2 ]);
	buf b_b_x_in_3 	(b_x_in[3 ], b_dinx[3 ]);
	buf b_b_x_in_4 	(b_x_in[4 ], b_dinx[4 ]);
	buf b_b_x_in_5 	(b_x_in[5 ], b_dinx[5 ]);
	buf b_b_x_in_6 	(b_x_in[6 ], b_dinx[6 ]);
	buf b_b_x_in_7 	(b_x_in[7 ], b_dinx[7 ]);
	buf b_b_x_in_8 	(b_x_in[8 ], b_dinx[8 ]);
	buf b_b_x_in_9 	(b_x_in[9 ], b_dinx[9 ]);
	buf b_b_x_in_10 (b_x_in[10], b_dinx[10]);
	buf b_b_x_in_11 (b_x_in[11], b_dinx[11]);	
	buf b_b_x_in_12 (b_x_in[12], b_dinx[12]);	
	  
	buf b_b_y_in_0 	(b_y_in[0 ], b_diny[0 ]);
	buf b_b_y_in_1 	(b_y_in[1 ], b_diny[1 ]);
	buf b_b_y_in_2 	(b_y_in[2 ], b_diny[2 ]);
	buf b_b_y_in_3 	(b_y_in[3 ], b_diny[3 ]);
	buf b_b_y_in_4 	(b_y_in[4 ], b_diny[4 ]);
	buf b_b_y_in_5 	(b_y_in[5 ], b_diny[5 ]);
	buf b_b_y_in_6 	(b_y_in[6 ], b_diny[6 ]);
	buf b_b_y_in_7 	(b_y_in[7 ], b_diny[7 ]);
	buf b_b_y_in_8 	(b_y_in[8 ], b_diny[8 ]);
	buf b_b_y_in_9 	(b_y_in[9 ], b_diny[9 ]);
	 
	buf b_b_z_in_0 	(b_z_in[0  ], b_dinz[0 ]);
	buf b_b_z_in_1 	(b_z_in[1  ], b_dinz[1 ]);
	buf b_b_z_in_2 	(b_z_in[2  ], b_dinz[2 ]);
	buf b_b_z_in_3 	(b_z_in[3  ], b_dinz[3 ]);
	buf b_b_z_in_4 	(b_z_in[4  ], b_dinz[4 ]);
	buf b_b_z_in_5 	(b_z_in[5  ], b_dinz[5 ]);
	buf b_b_z_in_6 	(b_z_in[6  ], b_dinz[6 ]);
	buf b_b_z_in_7 	(b_z_in[7  ], b_dinz[7 ]);
	buf b_b_z_in_8 	(b_z_in[8  ], b_dinz[8 ]);
	buf b_b_z_in_9 	(b_z_in[9  ], b_dinz[9 ]);
	buf b_b_z_in_10 (b_z_in[10 ], b_dinz[10]);
	buf b_b_z_in_11 (b_z_in[11 ], b_dinz[11]);	
	buf b_b_z_in_12 (b_z_in[12 ], b_dinz[12]);
	buf b_b_z_in_13 (b_z_in[13 ], b_dinz[13]);
	buf b_b_z_in_14 (b_z_in[14 ], b_dinz[14]);
	buf b_b_z_in_15 (b_z_in[15 ], b_dinz[15]);
	buf b_b_z_in_16 (b_z_in[16 ], b_dinz[16]);
	buf b_b_z_in_17 (b_z_in[17 ], b_dinz[17]);
	buf b_b_z_in_18 (b_z_in[18 ], b_dinz[18]);
	buf b_b_z_in_19 (b_z_in[19 ], b_dinz[19]);
	buf b_b_z_in_20 (b_z_in[20 ], b_dinz[20]);
	buf b_b_z_in_21 (b_z_in[21 ], b_dinz[21]);
	buf b_b_z_in_22 (b_z_in[22 ], b_dinz[22]);
	buf b_b_z_in_23 (b_z_in[23 ], b_dinz[23]);
	buf b_b_z_in_24 (b_z_in[24 ], b_dinz[24]);
	
	buf b_a_mac_out0  (a_mac_out[0  ], a_mac_o_out[0 ]);
	buf b_a_mac_out1  (a_mac_out[1  ], a_mac_o_out[1 ]);
	buf b_a_mac_out2  (a_mac_out[2  ], a_mac_o_out[2 ]);
	buf b_a_mac_out3  (a_mac_out[3  ], a_mac_o_out[3 ]);
	buf b_a_mac_out4  (a_mac_out[4  ], a_mac_o_out[4 ]);
	buf b_a_mac_out5  (a_mac_out[5  ], a_mac_o_out[5 ]);
	buf b_a_mac_out6  (a_mac_out[6  ], a_mac_o_out[6 ]);
	buf b_a_mac_out7  (a_mac_out[7  ], a_mac_o_out[7 ]);
	buf b_a_mac_out8  (a_mac_out[8  ], a_mac_o_out[8 ]);
	buf b_a_mac_out9  (a_mac_out[9  ], a_mac_o_out[9 ]);
	buf b_a_mac_out10 (a_mac_out[10 ], a_mac_o_out[10]);
	buf b_a_mac_out11 (a_mac_out[11 ], a_mac_o_out[11]);
	buf b_a_mac_out12 (a_mac_out[12 ], a_mac_o_out[12]);
	buf b_a_mac_out13 (a_mac_out[13 ], a_mac_o_out[13]);
	buf b_a_mac_out14 (a_mac_out[14 ], a_mac_o_out[14]);
	buf b_a_mac_out15 (a_mac_out[15 ], a_mac_o_out[15]);
	buf b_a_mac_out16 (a_mac_out[16 ], a_mac_o_out[16]);
	buf b_a_mac_out17 (a_mac_out[17 ], a_mac_o_out[17]);
	buf b_a_mac_out18 (a_mac_out[18 ], a_mac_o_out[18]);
	buf b_a_mac_out19 (a_mac_out[19 ], a_mac_o_out[19]);
	buf b_a_mac_out20 (a_mac_out[20 ], a_mac_o_out[20]);
	buf b_a_mac_out21 (a_mac_out[21 ], a_mac_o_out[21]);
	buf b_a_mac_out22 (a_mac_out[22 ], a_mac_o_out[22]);
	buf b_a_mac_out23 (a_mac_out[23 ], a_mac_o_out[23]);
	buf b_a_mac_out24 (a_mac_out[24 ], a_mac_o_out[24]);
	
	buf b_b_mac_out0  (b_mac_out[0  ], b_mac_o_out[0 ]);
	buf b_b_mac_out1  (b_mac_out[1  ], b_mac_o_out[1 ]);
	buf b_b_mac_out2  (b_mac_out[2  ], b_mac_o_out[2 ]);
	buf b_b_mac_out3  (b_mac_out[3  ], b_mac_o_out[3 ]);
	buf b_b_mac_out4  (b_mac_out[4  ], b_mac_o_out[4 ]);
	buf b_b_mac_out5  (b_mac_out[5  ], b_mac_o_out[5 ]);
	buf b_b_mac_out6  (b_mac_out[6  ], b_mac_o_out[6 ]);
	buf b_b_mac_out7  (b_mac_out[7  ], b_mac_o_out[7 ]);
	buf b_b_mac_out8  (b_mac_out[8  ], b_mac_o_out[8 ]);
	buf b_b_mac_out9  (b_mac_out[9  ], b_mac_o_out[9 ]);
	buf b_b_mac_out10 (b_mac_out[10 ], b_mac_o_out[10]);
	buf b_b_mac_out11 (b_mac_out[11 ], b_mac_o_out[11]);
	buf b_b_mac_out12 (b_mac_out[12 ], b_mac_o_out[12]);
	buf b_b_mac_out13 (b_mac_out[13 ], b_mac_o_out[13]);
	buf b_b_mac_out14 (b_mac_out[14 ], b_mac_o_out[14]);
	buf b_b_mac_out15 (b_mac_out[15 ], b_mac_o_out[15]);
	buf b_b_mac_out16 (b_mac_out[16 ], b_mac_o_out[16]);
	buf b_b_mac_out17 (b_mac_out[17 ], b_mac_o_out[17]);
	buf b_b_mac_out18 (b_mac_out[18 ], b_mac_o_out[18]);
	buf b_b_mac_out19 (b_mac_out[19 ], b_mac_o_out[19]);
	buf b_b_mac_out20 (b_mac_out[20 ], b_mac_o_out[20]);
	buf b_b_mac_out21 (b_mac_out[21 ], b_mac_o_out[21]);
	buf b_b_mac_out22 (b_mac_out[22 ], b_mac_o_out[22]);
	buf b_b_mac_out23 (b_mac_out[23 ], b_mac_o_out[23]);
	buf b_b_mac_out24 (b_mac_out[24 ], b_mac_o_out[24]);
	
	buf b_a_sload (a_sload_i, a_sload);
	buf b_a_acc_en (a_acc_en_i, a_acc_en);
	//buf b_a_dinz_en (a_dinz_en_i, a_dinz_en);
	
	buf b_b_sload   (b_sload_i,   b_sload);
	buf b_b_acc_en  (b_acc_en_i,  b_acc_en);
	//buf b_b_dinz_en (b_dinz_en_i, b_dinz_en);	   
    
	//*** Input a register x with 1 level deep of register

	always @(posedge clk_in or negedge a_in_rstn or negedge a_in_setn) begin
		if (!a_in_rstn)
			a_qx_o_reg_asyn <= 13'b0;
		else if(!a_in_setn)
			a_qx_o_reg_asyn <= 13'h1FFF;
		else if(a_dinxy_cen)
			a_qx_o_reg_asyn <= a_x_in;
	end

	always @(posedge clk_in) begin
		if (!a_in_rstn)
			a_qx_o_reg_syn <= 13'b0;
		else if(!a_in_setn)
			a_qx_o_reg_syn <= 13'h1FFF;
		else if(a_dinxy_cen)
			a_qx_o_reg_syn <= a_x_in;
	end
	assign a_qx_o_reg = a_sr_syn_sel == 1'b1 ? a_qx_o_reg_syn : a_qx_o_reg_asyn ;

	always @(a_x_in or a_qx_o_reg or a_xreg) begin
		case (a_xreg)
  	                0 : a_qx_o_mux <= a_x_in;
  	                1 : a_qx_o_mux <= a_qx_o_reg;
		endcase
	end

	//*** Input a register y with 1 level deep of registers
	always @(posedge clk_in or negedge a_in_rstn or negedge a_in_setn) begin
		if (!a_in_rstn)
			a_qy_o_reg_asyn <= 10'b0;
		else if(!a_in_setn)
			a_qy_o_reg_asyn <= 10'h3FF;
		else if(a_dinxy_cen)
			a_qy_o_reg_asyn <= a_y_in;
	end

	always @(posedge clk_in) begin
		if (!a_in_rstn)
			a_qy_o_reg_syn <= 10'b0;
		else if(!a_in_setn)
			a_qy_o_reg_syn <= 10'h3FF;
		else if(a_dinxy_cen)
			a_qy_o_reg_syn <= a_y_in;
	end
	assign a_qy_o_reg = a_sr_syn_sel == 1'b1 ? a_qy_o_reg_syn : a_qy_o_reg_asyn;

	always @(a_y_in or a_qy_o_reg or a_yreg) begin
		case (a_yreg)
  	                0 : a_qy_o_mux <= a_y_in;
  	                1 : a_qy_o_mux <= a_qy_o_reg;
		endcase
	end

	//*** Input a register z with 1 level deep of registers

	always @(posedge clk_in or negedge a_in_rstn or negedge a_in_setn) begin
		if (!a_in_rstn)
			a_qz_o_reg_asyn <= 25'b0;
		else if(!a_in_setn)
			a_qz_o_reg_asyn <= 25'h1FF_FFFF;
		else if(a_dinz_cen)
			a_qz_o_reg_asyn <= a_z_in;
	end

	always @(posedge clk_in) begin
		if (!a_in_rstn)
			a_qz_o_reg_syn <= 25'b0;
		else if(!a_in_setn)
			a_qz_o_reg_syn <= 25'h1FF_FFFF;
		else if(a_dinz_cen)
			a_qz_o_reg_syn <= a_z_in;
	end
	assign a_qz_o_reg = a_sr_syn_sel == 1'b1 ? a_qz_o_reg_syn : a_qz_o_reg_asyn ;

	always @(a_z_in or a_qz_o_reg or a_zreg) begin
		case (a_zreg)
  	                0 : a_qz_o_mux <= a_z_in;
  	                1 : a_qz_o_mux <= a_qz_o_reg;
		endcase
	end


	always @(posedge clk_in or negedge a_in_rstn) begin
		if (!a_in_rstn)
			a_dinz_en_reg_asyn <= 1'b0;
		else 
			a_dinz_en_reg_asyn <= a_dinz_en;
	end

	always @(posedge clk_in) begin
		if (!a_in_rstn)
			a_dinz_en_reg_syn <= 1'b0;
		else 
			a_dinz_en_reg_syn <= a_dinz_en;
	end
	assign a_dinz_en_reg = a_sr_syn_sel == 1'b1 ? a_dinz_en_reg_syn : a_dinz_en_reg_asyn ;

	always @(a_dinz_en or a_dinz_en_reg or a_zreg) begin
		case (a_zreg)
  	                0 : a_dinz_en_i <= a_dinz_en;
  	                1 : a_dinz_en_i <= a_dinz_en_reg;
		endcase
	end

	/*mac a	*/	
	//*** 12x9 Multiplier
	assign a_mult_o = (modea_sel == "12x9" || modea_sel == 3'b010)?{{12{a_signedx}}, a_qx_o_mux} * {{15{a_signedy}}, a_qy_o_mux}:0;

	//*** 25+25 adder
	assign a_add_o = (modea_sel == "12x9" || modea_sel == 3'b010)?((a_sload_i==1)?a_add_mux:(a_mult_o + a_add_mux)):0;

	//*** generate a_overflow
	assign a_overflow_tmp = (~(a_mult_o[24] ^ a_add_mux[24])) && (a_add_o[24] ^ a_add_mux[24]);

	always @(posedge clk_in or negedge a_ovf_rstn) begin
		if (!a_ovf_rstn)
  	          mac_a_overflow_d_asyn <= 1'b0;
		else if(a_mac_out_cen & mac_a_overflow_d_asyn)
  	          mac_a_overflow_d_asyn <= 1'b1;
		else if(a_mac_out_cen == 1'b0)
			  mac_a_overflow_d_asyn <= mac_a_overflow_d_asyn ;
		else
			  mac_a_overflow_d_asyn <= a_overflow_tmp ;
	end

	always @(posedge clk_in) begin
		if (!a_ovf_rstn)
  	          mac_a_overflow_d_syn <= 1'b0;
		else if(a_mac_out_cen & mac_a_overflow_d_syn)
  	          mac_a_overflow_d_syn <= 1'b1;
		else if(a_mac_out_cen == 1'b0)
			  mac_a_overflow_d_syn <= mac_a_overflow_d_syn ;	  
		else
			  mac_a_overflow_d_syn <= a_overflow_tmp ;
	end
	assign mac_a_overflow_d = a_sr_syn_sel == 1 ? mac_a_overflow_d_syn :  mac_a_overflow_d_asyn;

	always @(posedge clk_in or negedge a_out_sr) begin
		if (!a_out_sr)
  	          mac_a_overflow_temp_asyn <= 1'b0;
		else if(a_overflow_tmp)
  	          mac_a_overflow_temp_asyn <= 1'b1;
	end
	assign mac_a_overflow_or = mac_a_overflow_temp_asyn | a_overflow_tmp ;


    assign mac_a_overflow = a_macreg ? mac_a_overflow_d : mac_a_overflow_or;
    

	//*** adder/acc with 1 level of register
	mac_dff_sync dff_sync_a_0 (   .q(a_qmac_o_reg_syn[0]),.clk(clk_in),.d(a_qmac_i[0]),.rstn(a_6_out_rstn), .setn(a_6_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_1 (   .q(a_qmac_o_reg_syn[1]),.clk(clk_in),.d(a_qmac_i[1]),.rstn(a_7_out_rstn), .setn(a_7_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_2 (   .q(a_qmac_o_reg_syn[2]),.clk(clk_in),.d(a_qmac_i[2]),.rstn(a_8_out_rstn), .setn(a_8_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_3 (   .q(a_qmac_o_reg_syn[3]),.clk(clk_in),.d(a_qmac_i[3]),.rstn(a_9_out_rstn), .setn(a_9_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_4 (   .q(a_qmac_o_reg_syn[4]),.clk(clk_in),.d(a_qmac_i[4]),.rstn(a_10_out_rstn),.setn(a_10_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_5 (   .q(a_qmac_o_reg_syn[5]),.clk(clk_in),.d(a_qmac_i[5]),.rstn(a_11_out_rstn),.setn(a_11_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_6 (   .q(a_qmac_o_reg_syn[6]),.clk(clk_in),.d(a_qmac_i[6]),.rstn(a_12_out_rstn),.setn(a_12_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_7 (   .q(a_qmac_o_reg_syn[7]),.clk(clk_in),.d(a_qmac_i[7]),.rstn(a_13_out_rstn),.setn(a_13_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_8 (   .q(a_qmac_o_reg_syn[8]),.clk(clk_in),.d(a_qmac_i[8]),.rstn(a_14_out_rstn),.setn(a_14_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_9 (   .q(a_qmac_o_reg_syn[9]),.clk(clk_in),.d(a_qmac_i[9]),.rstn(a_15_out_rstn),.setn(a_15_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_10 (.q(a_qmac_o_reg_syn[10]),.clk(clk_in),.d(a_qmac_i[10]),.rstn(a_16_out_rstn),.setn(a_16_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_11 (.q(a_qmac_o_reg_syn[11]),.clk(clk_in),.d(a_qmac_i[11]),.rstn(a_17_out_rstn),.setn(a_17_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_12 (.q(a_qmac_o_reg_syn[12]),.clk(clk_in),.d(a_qmac_i[12]),.rstn(a_18_out_rstn),.setn(a_18_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_13 (.q(a_qmac_o_reg_syn[13]),.clk(clk_in),.d(a_qmac_i[13]),.rstn(a_19_out_rstn),.setn(a_19_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_14 (.q(a_qmac_o_reg_syn[14]),.clk(clk_in),.d(a_qmac_i[14]),.rstn(a_20_out_rstn),.setn(a_20_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_15 (.q(a_qmac_o_reg_syn[15]),.clk(clk_in),.d(a_qmac_i[15]),.rstn(a_21_out_rstn),.setn(a_21_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_16 (.q(a_qmac_o_reg_syn[16]),.clk(clk_in),.d(a_qmac_i[16]),.rstn(a_22_out_rstn),.setn(a_22_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_17 (.q(a_qmac_o_reg_syn[17]),.clk(clk_in),.d(a_qmac_i[17]),.rstn(a_23_out_rstn),.setn(a_23_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_18 (.q(a_qmac_o_reg_syn[18]),.clk(clk_in),.d(a_qmac_i[18]),.rstn(a_24_out_rstn),.setn(a_24_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_19 (.q(a_qmac_o_reg_syn[19]),.clk(clk_in),.d(a_qmac_i[19]),.rstn(a_25_out_rstn),.setn(a_25_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_20 (.q(a_qmac_o_reg_syn[20]),.clk(clk_in),.d(a_qmac_i[20]),.rstn(a_26_out_rstn),.setn(a_26_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_21 (.q(a_qmac_o_reg_syn[21]),.clk(clk_in),.d(a_qmac_i[21]),.rstn(a_27_out_rstn),.setn(a_27_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_22 (.q(a_qmac_o_reg_syn[22]),.clk(clk_in),.d(a_qmac_i[22]),.rstn(a_28_out_rstn),.setn(a_28_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_23 (.q(a_qmac_o_reg_syn[23]),.clk(clk_in),.d(a_qmac_i[23]),.rstn(a_29_out_rstn),.setn(a_29_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_a_24 (.q(a_qmac_o_reg_syn[24]),.clk(clk_in),.d(a_qmac_i[24]),.rstn(a_30_out_rstn),.setn(a_30_out_setn),.cen(a_mac_out_cen));

	mac_dff_async dff_async_a_0 (   .q(a_qmac_o_reg_asyn[0]),.clk(clk_in),.d(a_qmac_i[0]),.rstn(a_6_out_rstn), .setn(a_6_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_1 (   .q(a_qmac_o_reg_asyn[1]),.clk(clk_in),.d(a_qmac_i[1]),.rstn(a_7_out_rstn), .setn(a_7_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_2 (   .q(a_qmac_o_reg_asyn[2]),.clk(clk_in),.d(a_qmac_i[2]),.rstn(a_8_out_rstn), .setn(a_8_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_3 (   .q(a_qmac_o_reg_asyn[3]),.clk(clk_in),.d(a_qmac_i[3]),.rstn(a_9_out_rstn), .setn(a_9_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_4 (   .q(a_qmac_o_reg_asyn[4]),.clk(clk_in),.d(a_qmac_i[4]),.rstn(a_10_out_rstn),.setn(a_10_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_5 (   .q(a_qmac_o_reg_asyn[5]),.clk(clk_in),.d(a_qmac_i[5]),.rstn(a_11_out_rstn),.setn(a_11_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_6 (   .q(a_qmac_o_reg_asyn[6]),.clk(clk_in),.d(a_qmac_i[6]),.rstn(a_12_out_rstn),.setn(a_12_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_7 (   .q(a_qmac_o_reg_asyn[7]),.clk(clk_in),.d(a_qmac_i[7]),.rstn(a_13_out_rstn),.setn(a_13_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_8 (   .q(a_qmac_o_reg_asyn[8]),.clk(clk_in),.d(a_qmac_i[8]),.rstn(a_14_out_rstn),.setn(a_14_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_9 (   .q(a_qmac_o_reg_asyn[9]),.clk(clk_in),.d(a_qmac_i[9]),.rstn(a_15_out_rstn),.setn(a_15_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_10 (.q(a_qmac_o_reg_asyn[10]),.clk(clk_in),.d(a_qmac_i[10]),.rstn(a_16_out_rstn),.setn(a_16_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_11 (.q(a_qmac_o_reg_asyn[11]),.clk(clk_in),.d(a_qmac_i[11]),.rstn(a_17_out_rstn),.setn(a_17_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_12 (.q(a_qmac_o_reg_asyn[12]),.clk(clk_in),.d(a_qmac_i[12]),.rstn(a_18_out_rstn),.setn(a_18_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_13 (.q(a_qmac_o_reg_asyn[13]),.clk(clk_in),.d(a_qmac_i[13]),.rstn(a_19_out_rstn),.setn(a_19_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_14 (.q(a_qmac_o_reg_asyn[14]),.clk(clk_in),.d(a_qmac_i[14]),.rstn(a_20_out_rstn),.setn(a_20_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_15 (.q(a_qmac_o_reg_asyn[15]),.clk(clk_in),.d(a_qmac_i[15]),.rstn(a_21_out_rstn),.setn(a_21_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_16 (.q(a_qmac_o_reg_asyn[16]),.clk(clk_in),.d(a_qmac_i[16]),.rstn(a_22_out_rstn),.setn(a_22_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_17 (.q(a_qmac_o_reg_asyn[17]),.clk(clk_in),.d(a_qmac_i[17]),.rstn(a_23_out_rstn),.setn(a_23_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_18 (.q(a_qmac_o_reg_asyn[18]),.clk(clk_in),.d(a_qmac_i[18]),.rstn(a_24_out_rstn),.setn(a_24_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_19 (.q(a_qmac_o_reg_asyn[19]),.clk(clk_in),.d(a_qmac_i[19]),.rstn(a_25_out_rstn),.setn(a_25_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_20 (.q(a_qmac_o_reg_asyn[20]),.clk(clk_in),.d(a_qmac_i[20]),.rstn(a_26_out_rstn),.setn(a_26_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_21 (.q(a_qmac_o_reg_asyn[21]),.clk(clk_in),.d(a_qmac_i[21]),.rstn(a_27_out_rstn),.setn(a_27_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_22 (.q(a_qmac_o_reg_asyn[22]),.clk(clk_in),.d(a_qmac_i[22]),.rstn(a_28_out_rstn),.setn(a_28_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_23 (.q(a_qmac_o_reg_asyn[23]),.clk(clk_in),.d(a_qmac_i[23]),.rstn(a_29_out_rstn),.setn(a_29_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_a_24 (.q(a_qmac_o_reg_asyn[24]),.clk(clk_in),.d(a_qmac_i[24]),.rstn(a_30_out_rstn),.setn(a_30_out_setn),.cen(a_mac_out_cen));

	assign a_qmac_i = a_add_o ;
	assign a_qmac_o_reg = a_sr_syn_sel == 1 ? a_qmac_o_reg_syn :  a_qmac_o_reg_asyn ;
	always @(a_acc_en_i or a_dinz_en_i or a_qz_o_mux or a_qmac_o_reg or a_sload_i) begin
		if(a_sload_i == 1'b1)
			a_add_mux = a_qz_o_mux ;
		else if(a_acc_en_i == 1'b1)
			a_add_mux = a_qmac_o_reg ;
		else if(a_dinz_en_i == 1'b1)
			a_add_mux = a_qz_o_mux ;
		else
			a_add_mux = 25'b0;
	end

	
	//*** a mac output
	assign a_mac_o_mux = (modea_sel == "12x9" || modea_sel == 3'b010)?a_macreg?a_qmac_o_reg:a_add_o:0;	

	/*mac a	*/	
	
	//*** Input b register x with 1 level deep of register

	always @(posedge clk_in or negedge b_in_rstn or negedge b_in_setn) begin
		if (!b_in_rstn)
			b_qx_o_reg_asyn <= 13'b0;
		else if(!b_in_setn)
			b_qx_o_reg_asyn <= 13'h1FFF;
		else if(b_dinxy_cen)
			b_qx_o_reg_asyn <= b_x_in;
	end

	always @(posedge clk_in) begin
		if (!b_in_rstn)
			b_qx_o_reg_syn <= 13'b0;
		else if(!b_in_setn)
			b_qx_o_reg_syn <= 13'h1FFF;
		else if(b_dinxy_cen)
			b_qx_o_reg_syn <= b_x_in;
	end
	assign b_qx_o_reg = b_sr_syn_sel == 1 ? b_qx_o_reg_syn : b_qx_o_reg_asyn ;

	always @(b_x_in or b_qx_o_reg or b_xreg) begin
		case (b_xreg)
  	                0 : b_qx_o_mux <= b_x_in;
  	                1 : b_qx_o_mux <= b_qx_o_reg;
		endcase
	end

	//*** Input b register y with 1 level deep of registers

	always @(posedge clk_in or negedge b_in_rstn or negedge b_in_setn) begin
		if (!b_in_rstn)
			b_qy_o_reg_asyn <= 10'b0;
		else if(!b_in_setn)
			b_qy_o_reg_asyn <= 10'h3FF;
		else if(b_dinxy_cen)
			b_qy_o_reg_asyn <= b_y_in;
	end

	always @(posedge clk_in) begin
		if (!b_in_rstn)
			b_qy_o_reg_syn <= 10'b0;
		else if(!b_in_setn)
			b_qy_o_reg_syn <= 10'h3FF;
		else if(b_dinxy_cen)
			b_qy_o_reg_syn <= b_y_in;
	end
	assign b_qy_o_reg = b_sr_syn_sel == 1 ? b_qy_o_reg_syn : b_qy_o_reg_asyn ;
	always @(b_y_in or b_qy_o_reg or b_yreg) begin
		case (b_yreg)
  	                0 : b_qy_o_mux <= b_y_in;
  	                1 : b_qy_o_mux <= b_qy_o_reg;
		endcase
	end

	//*** Input b register z with 1 level deep of registers

	always @(posedge clk_in or negedge b_in_rstn or negedge b_in_setn) begin
		if (!b_in_rstn)
			b_qz_o_reg_asyn <= 25'b0;
		else if(!b_in_setn)
			b_qz_o_reg_asyn <= 25'h1FF_FFFF;
		else if(b_dinz_cen)
			b_qz_o_reg_asyn <= b_z_in;
	end

	always @(posedge clk_in) begin
		if (!b_in_rstn)
			b_qz_o_reg_syn <= 25'b0;
		else if(!b_in_setn)
			b_qz_o_reg_syn <= 25'h1FF_FFFF;
		else if(b_dinz_cen)
			b_qz_o_reg_syn <= b_z_in;
	end
	assign b_qz_o_reg = b_sr_syn_sel == 1 ? b_qz_o_reg_syn : b_qz_o_reg_asyn ;

	always @(b_z_in or b_qz_o_reg or b_zreg) begin
		case (b_zreg)
  	                0 : b_qz_o_mux <= b_z_in;
  	                1 : b_qz_o_mux <= b_qz_o_reg;
		endcase
	end


	always @(posedge clk_in or negedge b_in_rstn) begin
		if (!b_in_rstn)
			b_dinz_en_reg_asyn <= 1'b0;
		else 
			b_dinz_en_reg_asyn <= b_dinz_en;
	end

	always @(posedge clk_in) begin
		if (!b_in_rstn)
			b_dinz_en_reg_syn <= 1'b0;
		else 
			b_dinz_en_reg_syn <= b_dinz_en;
	end
	assign b_dinz_en_reg = b_sr_syn_sel == 1 ? b_dinz_en_reg_syn : b_dinz_en_reg_asyn ;

	always @(b_dinz_en or b_dinz_en_reg or b_zreg) begin
		case (b_zreg)
  	                0 : b_dinz_en_i <= b_dinz_en;
  	                1 : b_dinz_en_i <= b_dinz_en_reg;
		endcase
	end


	/*mac b	*/	
	//*** 12x9 Multiplier
	assign b_mult_o = (modeb_sel == "12x9" || modeb_sel == 3'b010)?{{12{b_signedx}}, b_qx_o_mux} * {{15{b_signedy}}, b_qy_o_mux}:0;

	//*** 25+25 adder
	assign b_add_o = (modeb_sel == "12x9" || modeb_sel == 3'b010)?((b_sload_i == 1)?b_add_mux:(b_mult_o + b_add_mux)):0;

	//*** generate b_overflow
	assign b_overflow_tmp = (~(b_mult_o[24] ^ b_add_mux[24])) && (b_add_o[24] ^ b_add_mux[24]);

	always @(posedge clk_in or negedge b_ovf_rstn) begin
		if (!b_ovf_rstn)
  	          mac_b_overflow_d_asyn <= 1'b0;
		else if(b_mac_out_cen & mac_b_overflow_d_asyn)
  	          mac_b_overflow_d_asyn <= 1'b1;
		else if(b_mac_out_cen == 1'b0)	  
			  mac_b_overflow_d_asyn <= mac_b_overflow_d_asyn ;
		else
			  mac_b_overflow_d_asyn <= b_overflow_tmp ;
	end

	always @(posedge clk_in) begin
		if (!b_ovf_rstn)
  	          mac_b_overflow_d_syn <= 1'b0;
		else if(b_mac_out_cen & mac_b_overflow_d_syn)
  	          mac_b_overflow_d_syn <= 1'b1;
		else if(b_mac_out_cen == 1'b0)	  
			  mac_b_overflow_d_syn <= mac_b_overflow_d_syn ;
		else
			  mac_b_overflow_d_syn <= b_overflow_tmp ;
	end
	assign mac_b_overflow_d = b_sr_syn_sel == 1 ? mac_b_overflow_d_syn : mac_b_overflow_d_asyn ;
	
	always @(posedge clk_in or negedge b_out_sr) begin
		if (!b_out_sr)
  	          mac_b_overflow_temp_asyn <= 1'b0;
		else if(b_overflow_tmp)
  	          mac_b_overflow_temp_asyn <= 1'b1;
	end
	assign mac_b_overflow_or = mac_b_overflow_temp_asyn | b_overflow_tmp ;

    assign b_overflow = b_macreg ? mac_b_overflow_d : mac_b_overflow_or;


	//*** adder/acc with 1 level of register
	mac_dff_sync dff_sync_b_0 (.q(b_qmac_o_reg_syn[0]),.clk(clk_in),.d(b_qmac_i[0]),.rstn(b_0_out_rstn),.setn(b_0_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_1 (.q(b_qmac_o_reg_syn[1]),.clk(clk_in),.d(b_qmac_i[1]),.rstn(b_1_out_rstn),.setn(b_1_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_2 (.q(b_qmac_o_reg_syn[2]),.clk(clk_in),.d(b_qmac_i[2]),.rstn(b_2_out_rstn),.setn(b_2_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_3 (.q(b_qmac_o_reg_syn[3]),.clk(clk_in),.d(b_qmac_i[3]),.rstn(b_3_out_rstn),.setn(b_3_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_4 (.q(b_qmac_o_reg_syn[4]),.clk(clk_in),.d(b_qmac_i[4]),.rstn(b_4_out_rstn),.setn(b_4_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_5 (.q(b_qmac_o_reg_syn[5]),.clk(clk_in),.d(b_qmac_i[5]),.rstn(b_5_out_rstn),.setn(b_5_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_6 (.q(b_qmac_o_reg_syn[6]),.clk(clk_in),.d(b_qmac_i[6]),.rstn(b_6_out_rstn),.setn(b_6_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_7 (.q(b_qmac_o_reg_syn[7]),.clk(clk_in),.d(b_qmac_i[7]),.rstn(b_7_out_rstn),.setn(b_7_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_8 (.q(b_qmac_o_reg_syn[8]),.clk(clk_in),.d(b_qmac_i[8]),.rstn(b_8_out_rstn),.setn(b_8_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_9 (.q(b_qmac_o_reg_syn[9]),.clk(clk_in),.d(b_qmac_i[9]),.rstn(b_9_out_rstn),.setn(b_9_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_10 (.q(b_qmac_o_reg_syn[10]),.clk(clk_in),.d(b_qmac_i[10]),.rstn(b_10_out_rstn),.setn(b_10_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_11 (.q(b_qmac_o_reg_syn[11]),.clk(clk_in),.d(b_qmac_i[11]),.rstn(b_11_out_rstn),.setn(b_11_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_12 (.q(b_qmac_o_reg_syn[12]),.clk(clk_in),.d(b_qmac_i[12]),.rstn(b_12_out_rstn),.setn(b_12_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_13 (.q(b_qmac_o_reg_syn[13]),.clk(clk_in),.d(b_qmac_i[13]),.rstn(b_13_out_rstn),.setn(b_13_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_14 (.q(b_qmac_o_reg_syn[14]),.clk(clk_in),.d(b_qmac_i[14]),.rstn(b_14_out_rstn),.setn(b_14_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_15 (.q(b_qmac_o_reg_syn[15]),.clk(clk_in),.d(b_qmac_i[15]),.rstn(b_15_out_rstn),.setn(b_15_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_16 (.q(b_qmac_o_reg_syn[16]),.clk(clk_in),.d(b_qmac_i[16]),.rstn(b_16_out_rstn),.setn(b_16_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_17 (.q(b_qmac_o_reg_syn[17]),.clk(clk_in),.d(b_qmac_i[17]),.rstn(b_17_out_rstn),.setn(b_17_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_18 (.q(b_qmac_o_reg_syn[18]),.clk(clk_in),.d(b_qmac_i[18]),.rstn(b_18_out_rstn),.setn(b_18_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_19 (.q(b_qmac_o_reg_syn[19]),.clk(clk_in),.d(b_qmac_i[19]),.rstn(b_19_out_rstn),.setn(b_19_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_20 (.q(b_qmac_o_reg_syn[20]),.clk(clk_in),.d(b_qmac_i[20]),.rstn(b_20_out_rstn),.setn(b_20_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_21 (.q(b_qmac_o_reg_syn[21]),.clk(clk_in),.d(b_qmac_i[21]),.rstn(b_21_out_rstn),.setn(b_21_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_22 (.q(b_qmac_o_reg_syn[22]),.clk(clk_in),.d(b_qmac_i[22]),.rstn(b_22_out_rstn),.setn(b_22_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_23 (.q(b_qmac_o_reg_syn[23]),.clk(clk_in),.d(b_qmac_i[23]),.rstn(b_23_out_rstn),.setn(b_23_out_setn),.cen(b_mac_out_cen));
	mac_dff_sync dff_sync_b_24 (.q(b_qmac_o_reg_syn[24]),.clk(clk_in),.d(b_qmac_i[24]),.rstn(b_24_out_rstn),.setn(b_24_out_setn),.cen(b_mac_out_cen));

	mac_dff_async dff_async_b_0 (.q(b_qmac_o_reg_asyn[0]),.clk(clk_in),.d(b_qmac_i[0]),.rstn(b_0_out_rstn),.setn(b_0_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_1 (.q(b_qmac_o_reg_asyn[1]),.clk(clk_in),.d(b_qmac_i[1]),.rstn(b_1_out_rstn),.setn(b_1_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_2 (.q(b_qmac_o_reg_asyn[2]),.clk(clk_in),.d(b_qmac_i[2]),.rstn(b_2_out_rstn),.setn(b_2_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_3 (.q(b_qmac_o_reg_asyn[3]),.clk(clk_in),.d(b_qmac_i[3]),.rstn(b_3_out_rstn),.setn(b_3_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_4 (.q(b_qmac_o_reg_asyn[4]),.clk(clk_in),.d(b_qmac_i[4]),.rstn(b_4_out_rstn),.setn(b_4_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_5 (.q(b_qmac_o_reg_asyn[5]),.clk(clk_in),.d(b_qmac_i[5]),.rstn(b_5_out_rstn),.setn(b_5_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_6 (.q(b_qmac_o_reg_asyn[6]),.clk(clk_in),.d(b_qmac_i[6]),.rstn(b_6_out_rstn),.setn(b_6_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_7 (.q(b_qmac_o_reg_asyn[7]),.clk(clk_in),.d(b_qmac_i[7]),.rstn(b_7_out_rstn),.setn(b_7_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_8 (.q(b_qmac_o_reg_asyn[8]),.clk(clk_in),.d(b_qmac_i[8]),.rstn(b_8_out_rstn),.setn(b_8_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_9 (.q(b_qmac_o_reg_asyn[9]),.clk(clk_in),.d(b_qmac_i[9]),.rstn(b_9_out_rstn),.setn(b_9_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_10 (.q(b_qmac_o_reg_asyn[10]),.clk(clk_in),.d(b_qmac_i[10]),.rstn(b_10_out_rstn),.setn(b_10_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_11 (.q(b_qmac_o_reg_asyn[11]),.clk(clk_in),.d(b_qmac_i[11]),.rstn(b_11_out_rstn),.setn(b_11_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_12 (.q(b_qmac_o_reg_asyn[12]),.clk(clk_in),.d(b_qmac_i[12]),.rstn(b_12_out_rstn),.setn(b_12_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_13 (.q(b_qmac_o_reg_asyn[13]),.clk(clk_in),.d(b_qmac_i[13]),.rstn(b_13_out_rstn),.setn(b_13_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_14 (.q(b_qmac_o_reg_asyn[14]),.clk(clk_in),.d(b_qmac_i[14]),.rstn(b_14_out_rstn),.setn(b_14_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_15 (.q(b_qmac_o_reg_asyn[15]),.clk(clk_in),.d(b_qmac_i[15]),.rstn(b_15_out_rstn),.setn(b_15_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_16 (.q(b_qmac_o_reg_asyn[16]),.clk(clk_in),.d(b_qmac_i[16]),.rstn(b_16_out_rstn),.setn(b_16_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_17 (.q(b_qmac_o_reg_asyn[17]),.clk(clk_in),.d(b_qmac_i[17]),.rstn(b_17_out_rstn),.setn(b_17_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_18 (.q(b_qmac_o_reg_asyn[18]),.clk(clk_in),.d(b_qmac_i[18]),.rstn(b_18_out_rstn),.setn(b_18_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_19 (.q(b_qmac_o_reg_asyn[19]),.clk(clk_in),.d(b_qmac_i[19]),.rstn(b_19_out_rstn),.setn(b_19_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_20 (.q(b_qmac_o_reg_asyn[20]),.clk(clk_in),.d(b_qmac_i[20]),.rstn(b_20_out_rstn),.setn(b_20_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_21 (.q(b_qmac_o_reg_asyn[21]),.clk(clk_in),.d(b_qmac_i[21]),.rstn(b_21_out_rstn),.setn(b_21_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_22 (.q(b_qmac_o_reg_asyn[22]),.clk(clk_in),.d(b_qmac_i[22]),.rstn(b_22_out_rstn),.setn(b_22_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_23 (.q(b_qmac_o_reg_asyn[23]),.clk(clk_in),.d(b_qmac_i[23]),.rstn(b_23_out_rstn),.setn(b_23_out_setn),.cen(b_mac_out_cen));
	mac_dff_async dff_async_b_24 (.q(b_qmac_o_reg_asyn[24]),.clk(clk_in),.d(b_qmac_i[24]),.rstn(b_24_out_rstn),.setn(b_24_out_setn),.cen(b_mac_out_cen));


	assign b_qmac_i = b_add_o ;
	assign b_qmac_o_reg =  b_sr_syn_sel == 1 ? b_qmac_o_reg_syn : b_qmac_o_reg_asyn ;
	always @(b_acc_en_i or b_dinz_en_i or b_qz_o_mux or b_qmac_o_reg or b_sload_i) begin
		if(b_sload_i == 1'b1)
			b_add_mux = b_qz_o_mux ;
		else if(b_acc_en_i == 1'b1)
			b_add_mux = b_qmac_o_reg;
		else if(b_dinz_en_i == 1'b1)
			b_add_mux = b_qz_o_mux ;
		else
			b_add_mux <= 25'b0 ;
	end
	
	//*** b mac output
	assign b_mac_o_mux = (modeb_sel == "12x9" || modeb_sel == 3'b010)?b_macreg?b_qmac_o_reg:b_add_o:0;	

	/*mac b	*/	
	
	/*mac 18x18	*/	
	assign qx_o_mux = (modea_sel == "18x18" || modea_sel == 3'b001)?{b_qx_o_mux[12:0],a_qx_o_mux[5:0]}:19'b0;
	assign qy_o_mux = (modea_sel == "18x18" || modea_sel == 3'b001)?{b_qy_o_mux[9:0],a_qy_o_mux[8:0]}:19'b0;
	assign qz_o_mux = (modea_sel == "18x18" || modea_sel == 3'b001)?{b_qz_o_mux[23:0],a_qz_o_mux[23:0]}:48'b0;
	//*** 18x18 Multiplier
	assign mult_o = (modea_sel == "18x18" || modea_sel == 3'b001)?{{30{signedx}}, qx_o_mux} * {{30{signedy}}, qy_o_mux}:48'b0;

	//*** 48+48 adder
	assign add_o = (modea_sel == "18x18" || modea_sel == 3'b001)?((sload_i == 1)?add_mux:(mult_o + add_mux)):0;

	//*** generate mac_overflow for 18x18
	assign mac_overflow_tmp = (~(mult_o[47] ^ add_mux[47])) && (add_o[47] ^ add_mux[47]);

	always @(posedge clk_in or negedge a_ovf_rstn) begin
		if (!a_ovf_rstn)
  	          mac_overflow_d_asyn <= 1'b0;
		else if(a_mac_out_cen & mac_overflow_d_asyn)
  	          mac_overflow_d_asyn <= 1'b1;
		else if(a_mac_out_cen == 1'b0)
			  mac_overflow_d_asyn <= mac_overflow_d_asyn ;
		else
			  mac_overflow_d_asyn <= mac_overflow_tmp ;
	end

	always @(posedge clk_in) begin
		if (!a_ovf_rstn)
  	          mac_overflow_d_syn <= 1'b0;
		else if(a_mac_out_cen & mac_overflow_d_syn)
  	          mac_overflow_d_syn <= 1'b1;
		else if(a_mac_out_cen == 1'b0)
			  mac_overflow_d_syn <= mac_overflow_d_syn ;	  
		else
			  mac_overflow_d_syn <= mac_overflow_tmp ;
	end
	assign mac_overflow_d = a_sr_syn_sel == 1 ? mac_overflow_d_syn : mac_overflow_d_asyn ;

	always @(posedge clk_in or negedge a_out_sr) begin
		if (!a_out_sr)
  	          mac_overflow_temp_asyn <= 1'b0;
		else if(mac_overflow_tmp)
  	          mac_overflow_temp_asyn <= 1'b1;
	end
	assign mac_overflow_or =  mac_overflow_temp_asyn | mac_overflow_tmp ;

    assign mac_overflow = a_macreg ? mac_overflow_d : mac_overflow_or;

	//*** adder/acc with 1 level of register
	assign qmac_i = add_o ;
	mac_dff_sync dff_sync_ab_0 (.q(qmac_o_reg_syn[0]),.clk(clk_in),.d(qmac_i[0]),.rstn(a_0_out_rstn),.setn(a_0_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_1 (.q(qmac_o_reg_syn[1]),.clk(clk_in),.d(qmac_i[1]),.rstn(a_1_out_rstn),.setn(a_1_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_2 (.q(qmac_o_reg_syn[2]),.clk(clk_in),.d(qmac_i[2]),.rstn(a_2_out_rstn),.setn(a_2_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_3 (.q(qmac_o_reg_syn[3]),.clk(clk_in),.d(qmac_i[3]),.rstn(a_3_out_rstn),.setn(a_3_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_4 (.q(qmac_o_reg_syn[4]),.clk(clk_in),.d(qmac_i[4]),.rstn(a_4_out_rstn),.setn(a_4_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_5 (.q(qmac_o_reg_syn[5]),.clk(clk_in),.d(qmac_i[5]),.rstn(a_5_out_rstn),.setn(a_5_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_6 (.q(qmac_o_reg_syn[6]),.clk(clk_in),.d(qmac_i[6]),.rstn(a_6_out_rstn),.setn(a_6_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_7 (.q(qmac_o_reg_syn[7]),.clk(clk_in),.d(qmac_i[7]),.rstn(a_7_out_rstn),.setn(a_7_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_8 (.q(qmac_o_reg_syn[8]),.clk(clk_in),.d(qmac_i[8]),.rstn(a_8_out_rstn),.setn(a_8_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_9 (.q(qmac_o_reg_syn[9]),.clk(clk_in),.d(qmac_i[9]),.rstn(a_9_out_rstn),.setn(a_9_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_10 (.q(qmac_o_reg_syn[10]),.clk(clk_in),.d(qmac_i[10]),.rstn(a_10_out_rstn),.setn(a_10_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_11 (.q(qmac_o_reg_syn[11]),.clk(clk_in),.d(qmac_i[11]),.rstn(a_11_out_rstn),.setn(a_11_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_12 (.q(qmac_o_reg_syn[12]),.clk(clk_in),.d(qmac_i[12]),.rstn(a_12_out_rstn),.setn(a_12_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_13 (.q(qmac_o_reg_syn[13]),.clk(clk_in),.d(qmac_i[13]),.rstn(a_13_out_rstn),.setn(a_13_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_14 (.q(qmac_o_reg_syn[14]),.clk(clk_in),.d(qmac_i[14]),.rstn(a_14_out_rstn),.setn(a_14_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_15 (.q(qmac_o_reg_syn[15]),.clk(clk_in),.d(qmac_i[15]),.rstn(a_15_out_rstn),.setn(a_15_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_16 (.q(qmac_o_reg_syn[16]),.clk(clk_in),.d(qmac_i[16]),.rstn(a_16_out_rstn),.setn(a_16_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_17 (.q(qmac_o_reg_syn[17]),.clk(clk_in),.d(qmac_i[17]),.rstn(a_17_out_rstn),.setn(a_17_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_18 (.q(qmac_o_reg_syn[18]),.clk(clk_in),.d(qmac_i[18]),.rstn(a_18_out_rstn),.setn(a_18_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_19 (.q(qmac_o_reg_syn[19]),.clk(clk_in),.d(qmac_i[19]),.rstn(a_19_out_rstn),.setn(a_19_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_20 (.q(qmac_o_reg_syn[20]),.clk(clk_in),.d(qmac_i[20]),.rstn(a_20_out_rstn),.setn(a_20_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_21 (.q(qmac_o_reg_syn[21]),.clk(clk_in),.d(qmac_i[21]),.rstn(a_21_out_rstn),.setn(a_21_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_22 (.q(qmac_o_reg_syn[22]),.clk(clk_in),.d(qmac_i[22]),.rstn(a_22_out_rstn),.setn(a_22_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_23 (.q(qmac_o_reg_syn[23]),.clk(clk_in),.d(qmac_i[23]),.rstn(a_23_out_rstn),.setn(a_23_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_24 (.q(qmac_o_reg_syn[24]),.clk(clk_in),.d(qmac_i[24]),.rstn(a_24_out_rstn),.setn(a_24_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_25 (.q(qmac_o_reg_syn[25]),.clk(clk_in),.d(qmac_i[25]),.rstn(a_25_out_rstn),.setn(a_25_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_26 (.q(qmac_o_reg_syn[26]),.clk(clk_in),.d(qmac_i[26]),.rstn(a_26_out_rstn),.setn(a_26_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_27 (.q(qmac_o_reg_syn[27]),.clk(clk_in),.d(qmac_i[27]),.rstn(a_27_out_rstn),.setn(a_27_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_28 (.q(qmac_o_reg_syn[28]),.clk(clk_in),.d(qmac_i[28]),.rstn(a_28_out_rstn),.setn(a_28_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_29 (.q(qmac_o_reg_syn[29]),.clk(clk_in),.d(qmac_i[29]),.rstn(a_29_out_rstn),.setn(a_29_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_30 (.q(qmac_o_reg_syn[30]),.clk(clk_in),.d(qmac_i[30]),.rstn(a_30_out_rstn),.setn(a_30_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_31 (.q(qmac_o_reg_syn[31]),.clk(clk_in),.d(qmac_i[31]),.rstn(a_31_out_rstn),.setn(a_31_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_32 (.q(qmac_o_reg_syn[32]),.clk(clk_in),.d(qmac_i[32]),.rstn(a_32_out_rstn),.setn(a_32_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_33 (.q(qmac_o_reg_syn[33]),.clk(clk_in),.d(qmac_i[33]),.rstn(a_33_out_rstn),.setn(a_33_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_34 (.q(qmac_o_reg_syn[34]),.clk(clk_in),.d(qmac_i[34]),.rstn(a_34_out_rstn),.setn(a_34_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_35 (.q(qmac_o_reg_syn[35]),.clk(clk_in),.d(qmac_i[35]),.rstn(a_35_out_rstn),.setn(a_35_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_36 (.q(qmac_o_reg_syn[36]),.clk(clk_in),.d(qmac_i[36]),.rstn(a_36_out_rstn),.setn(a_36_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_37 (.q(qmac_o_reg_syn[37]),.clk(clk_in),.d(qmac_i[37]),.rstn(a_37_out_rstn),.setn(a_37_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_38 (.q(qmac_o_reg_syn[38]),.clk(clk_in),.d(qmac_i[38]),.rstn(a_38_out_rstn),.setn(a_38_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_39 (.q(qmac_o_reg_syn[39]),.clk(clk_in),.d(qmac_i[39]),.rstn(a_39_out_rstn),.setn(a_39_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_40 (.q(qmac_o_reg_syn[40]),.clk(clk_in),.d(qmac_i[40]),.rstn(a_40_out_rstn),.setn(a_40_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_41 (.q(qmac_o_reg_syn[41]),.clk(clk_in),.d(qmac_i[41]),.rstn(a_41_out_rstn),.setn(a_41_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_42 (.q(qmac_o_reg_syn[42]),.clk(clk_in),.d(qmac_i[42]),.rstn(a_42_out_rstn),.setn(a_42_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_43 (.q(qmac_o_reg_syn[43]),.clk(clk_in),.d(qmac_i[43]),.rstn(a_43_out_rstn),.setn(a_43_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_44 (.q(qmac_o_reg_syn[44]),.clk(clk_in),.d(qmac_i[44]),.rstn(a_44_out_rstn),.setn(a_44_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_45 (.q(qmac_o_reg_syn[45]),.clk(clk_in),.d(qmac_i[45]),.rstn(a_45_out_rstn),.setn(a_45_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_46 (.q(qmac_o_reg_syn[46]),.clk(clk_in),.d(qmac_i[46]),.rstn(a_46_out_rstn),.setn(a_46_out_setn),.cen(a_mac_out_cen));
	mac_dff_sync dff_sync_ab_47 (.q(qmac_o_reg_syn[47]),.clk(clk_in),.d(qmac_i[47]),.rstn(a_47_out_rstn),.setn(a_47_out_setn),.cen(a_mac_out_cen));

	mac_dff_async dff_async_ab_0 (.q(qmac_o_reg_asyn[0]),.clk(clk_in),.d(qmac_i[0]),.rstn(a_0_out_rstn),.setn(a_0_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_1 (.q(qmac_o_reg_asyn[1]),.clk(clk_in),.d(qmac_i[1]),.rstn(a_1_out_rstn),.setn(a_1_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_2 (.q(qmac_o_reg_asyn[2]),.clk(clk_in),.d(qmac_i[2]),.rstn(a_2_out_rstn),.setn(a_2_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_3 (.q(qmac_o_reg_asyn[3]),.clk(clk_in),.d(qmac_i[3]),.rstn(a_3_out_rstn),.setn(a_3_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_4 (.q(qmac_o_reg_asyn[4]),.clk(clk_in),.d(qmac_i[4]),.rstn(a_4_out_rstn),.setn(a_4_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_5 (.q(qmac_o_reg_asyn[5]),.clk(clk_in),.d(qmac_i[5]),.rstn(a_5_out_rstn),.setn(a_5_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_6 (.q(qmac_o_reg_asyn[6]),.clk(clk_in),.d(qmac_i[6]),.rstn(a_6_out_rstn),.setn(a_6_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_7 (.q(qmac_o_reg_asyn[7]),.clk(clk_in),.d(qmac_i[7]),.rstn(a_7_out_rstn),.setn(a_7_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_8 (.q(qmac_o_reg_asyn[8]),.clk(clk_in),.d(qmac_i[8]),.rstn(a_8_out_rstn),.setn(a_8_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_9 (.q(qmac_o_reg_asyn[9]),.clk(clk_in),.d(qmac_i[9]),.rstn(a_9_out_rstn),.setn(a_9_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_10 (.q(qmac_o_reg_asyn[10]),.clk(clk_in),.d(qmac_i[10]),.rstn(a_10_out_rstn),.setn(a_10_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_11 (.q(qmac_o_reg_asyn[11]),.clk(clk_in),.d(qmac_i[11]),.rstn(a_11_out_rstn),.setn(a_11_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_12 (.q(qmac_o_reg_asyn[12]),.clk(clk_in),.d(qmac_i[12]),.rstn(a_12_out_rstn),.setn(a_12_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_13 (.q(qmac_o_reg_asyn[13]),.clk(clk_in),.d(qmac_i[13]),.rstn(a_13_out_rstn),.setn(a_13_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_14 (.q(qmac_o_reg_asyn[14]),.clk(clk_in),.d(qmac_i[14]),.rstn(a_14_out_rstn),.setn(a_14_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_15 (.q(qmac_o_reg_asyn[15]),.clk(clk_in),.d(qmac_i[15]),.rstn(a_15_out_rstn),.setn(a_15_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_16 (.q(qmac_o_reg_asyn[16]),.clk(clk_in),.d(qmac_i[16]),.rstn(a_16_out_rstn),.setn(a_16_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_17 (.q(qmac_o_reg_asyn[17]),.clk(clk_in),.d(qmac_i[17]),.rstn(a_17_out_rstn),.setn(a_17_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_18 (.q(qmac_o_reg_asyn[18]),.clk(clk_in),.d(qmac_i[18]),.rstn(a_18_out_rstn),.setn(a_18_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_19 (.q(qmac_o_reg_asyn[19]),.clk(clk_in),.d(qmac_i[19]),.rstn(a_19_out_rstn),.setn(a_19_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_20 (.q(qmac_o_reg_asyn[20]),.clk(clk_in),.d(qmac_i[20]),.rstn(a_20_out_rstn),.setn(a_20_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_21 (.q(qmac_o_reg_asyn[21]),.clk(clk_in),.d(qmac_i[21]),.rstn(a_21_out_rstn),.setn(a_21_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_22 (.q(qmac_o_reg_asyn[22]),.clk(clk_in),.d(qmac_i[22]),.rstn(a_22_out_rstn),.setn(a_22_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_23 (.q(qmac_o_reg_asyn[23]),.clk(clk_in),.d(qmac_i[23]),.rstn(a_23_out_rstn),.setn(a_23_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_24 (.q(qmac_o_reg_asyn[24]),.clk(clk_in),.d(qmac_i[24]),.rstn(a_24_out_rstn),.setn(a_24_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_25 (.q(qmac_o_reg_asyn[25]),.clk(clk_in),.d(qmac_i[25]),.rstn(a_25_out_rstn),.setn(a_25_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_26 (.q(qmac_o_reg_asyn[26]),.clk(clk_in),.d(qmac_i[26]),.rstn(a_26_out_rstn),.setn(a_26_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_27 (.q(qmac_o_reg_asyn[27]),.clk(clk_in),.d(qmac_i[27]),.rstn(a_27_out_rstn),.setn(a_27_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_28 (.q(qmac_o_reg_asyn[28]),.clk(clk_in),.d(qmac_i[28]),.rstn(a_28_out_rstn),.setn(a_28_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_29 (.q(qmac_o_reg_asyn[29]),.clk(clk_in),.d(qmac_i[29]),.rstn(a_29_out_rstn),.setn(a_29_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_30 (.q(qmac_o_reg_asyn[30]),.clk(clk_in),.d(qmac_i[30]),.rstn(a_30_out_rstn),.setn(a_30_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_31 (.q(qmac_o_reg_asyn[31]),.clk(clk_in),.d(qmac_i[31]),.rstn(a_31_out_rstn),.setn(a_31_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_32 (.q(qmac_o_reg_asyn[32]),.clk(clk_in),.d(qmac_i[32]),.rstn(a_32_out_rstn),.setn(a_32_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_33 (.q(qmac_o_reg_asyn[33]),.clk(clk_in),.d(qmac_i[33]),.rstn(a_33_out_rstn),.setn(a_33_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_34 (.q(qmac_o_reg_asyn[34]),.clk(clk_in),.d(qmac_i[34]),.rstn(a_34_out_rstn),.setn(a_34_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_35 (.q(qmac_o_reg_asyn[35]),.clk(clk_in),.d(qmac_i[35]),.rstn(a_35_out_rstn),.setn(a_35_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_36 (.q(qmac_o_reg_asyn[36]),.clk(clk_in),.d(qmac_i[36]),.rstn(a_36_out_rstn),.setn(a_36_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_37 (.q(qmac_o_reg_asyn[37]),.clk(clk_in),.d(qmac_i[37]),.rstn(a_37_out_rstn),.setn(a_37_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_38 (.q(qmac_o_reg_asyn[38]),.clk(clk_in),.d(qmac_i[38]),.rstn(a_38_out_rstn),.setn(a_38_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_39 (.q(qmac_o_reg_asyn[39]),.clk(clk_in),.d(qmac_i[39]),.rstn(a_39_out_rstn),.setn(a_39_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_40 (.q(qmac_o_reg_asyn[40]),.clk(clk_in),.d(qmac_i[40]),.rstn(a_40_out_rstn),.setn(a_40_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_41 (.q(qmac_o_reg_asyn[41]),.clk(clk_in),.d(qmac_i[41]),.rstn(a_41_out_rstn),.setn(a_41_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_42 (.q(qmac_o_reg_asyn[42]),.clk(clk_in),.d(qmac_i[42]),.rstn(a_42_out_rstn),.setn(a_42_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_43 (.q(qmac_o_reg_asyn[43]),.clk(clk_in),.d(qmac_i[43]),.rstn(a_43_out_rstn),.setn(a_43_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_44 (.q(qmac_o_reg_asyn[44]),.clk(clk_in),.d(qmac_i[44]),.rstn(a_44_out_rstn),.setn(a_44_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_45 (.q(qmac_o_reg_asyn[45]),.clk(clk_in),.d(qmac_i[45]),.rstn(a_45_out_rstn),.setn(a_45_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_46 (.q(qmac_o_reg_asyn[46]),.clk(clk_in),.d(qmac_i[46]),.rstn(a_46_out_rstn),.setn(a_46_out_setn),.cen(a_mac_out_cen));
	mac_dff_async dff_async_ab_47 (.q(qmac_o_reg_asyn[47]),.clk(clk_in),.d(qmac_i[47]),.rstn(a_47_out_rstn),.setn(a_47_out_setn),.cen(a_mac_out_cen));

	assign qmac_o_reg = a_sr_syn_sel == 1 ? qmac_o_reg_syn : qmac_o_reg_asyn ;
	//always @(acc_en_i or dinz_en_i or qz_o_mux or qmac_o_reg) begin
	//	case ({acc_en_i,dinz_en_i})
    //              2'b01 : add_mux <= qz_o_mux;
    //              2'b10 : add_mux <= qmac_o_reg;
    //              default:add_mux <= 40'b0;
	//	endcase
	//end
	always @(acc_en_i or dinz_en_i or qz_o_mux or qmac_o_reg or sload_i) begin
		if(sload_i == 1'b1)
			add_mux = qz_o_mux ;
		else if(acc_en_i)
			add_mux = qmac_o_reg ;
		else if(dinz_en_i)
			add_mux = qz_o_mux ;
		else
			add_mux = 48'b0;
	end
	
	//*** mac output
	assign mac_o_mux = (modea_sel == "18x18" || modea_sel == 3'b001)?macreg?qmac_o_reg:add_o:48'b0;	

	/*mac*/		
	assign a_mac_o_out = 	(modea_sel == "18x18" || modea_sel == 3'b001)?mac_o_mux[23:0]:
				(modea_sel == "12x9" || modea_sel == 3'b010)?a_mac_o_mux:0;
	assign b_mac_o_out = 	(modeb_sel == "18x18" || modeb_sel == 3'b001)?mac_o_mux[47:24]:
				(modeb_sel == "12x9" || modeb_sel == 3'b010)?b_mac_o_mux:0;
		
	//*** make mac_a_overflow and mac_overflow together be a_overflow
	assign a_overflow =	(modea_sel == "18x18" || modea_sel == 3'b001)?mac_overflow:
				(modea_sel == "12x9" || modea_sel == 3'b010)?mac_a_overflow:0; 
	specify
	//iopath
(clk          =>   a_mac_out[0]      ) = (0,0);
(clk          =>   a_mac_out[1]      ) = (0,0);
(clk          =>   a_mac_out[2]      ) = (0,0);
(clk          =>   a_mac_out[3]      ) = (0,0);
(clk          =>   a_mac_out[4]      ) = (0,0);
(clk          =>   a_mac_out[5]      ) = (0,0);
(clk          =>   a_mac_out[6]      ) = (0,0);
(clk          =>   a_mac_out[7]      ) = (0,0);
(clk          =>   a_mac_out[8]      ) = (0,0);
(clk          =>   a_mac_out[9]      ) = (0,0);
(clk          =>   a_mac_out[10]     ) = (0,0);
(clk          =>   a_mac_out[11]     ) = (0,0);
(clk          =>   a_mac_out[12]     ) = (0,0);
(clk          =>   a_mac_out[13]     ) = (0,0);
(clk          =>   a_mac_out[14]     ) = (0,0);
(clk          =>   a_mac_out[15]     ) = (0,0);
(clk          =>   a_mac_out[16]     ) = (0,0);
(clk          =>   a_mac_out[17]     ) = (0,0);
(clk          =>   a_mac_out[18]     ) = (0,0);
(clk          =>   a_mac_out[19]     ) = (0,0);
(clk          =>   a_mac_out[20]     ) = (0,0);
(clk          =>   a_mac_out[21]     ) = (0,0);
(clk          =>   a_mac_out[22]     ) = (0,0);
(clk          =>   a_mac_out[23]     ) = (0,0);
(clk          =>   b_mac_out[0]      ) = (0,0);
(clk          =>   b_mac_out[1]      ) = (0,0);
(clk          =>   b_mac_out[2]      ) = (0,0);
(clk          =>   b_mac_out[3]      ) = (0,0);
(clk          =>   b_mac_out[4]      ) = (0,0);
(clk          =>   b_mac_out[5]      ) = (0,0);
(clk          =>   b_mac_out[6]      ) = (0,0);
(clk          =>   b_mac_out[7]      ) = (0,0);
(clk          =>   b_mac_out[8]      ) = (0,0);
(clk          =>   b_mac_out[9]      ) = (0,0);
(clk          =>   b_mac_out[10]     ) = (0,0);
(clk          =>   b_mac_out[11]     ) = (0,0);
(clk          =>   b_mac_out[12]     ) = (0,0);
(clk          =>   b_mac_out[13]     ) = (0,0);
(clk          =>   b_mac_out[14]     ) = (0,0);
(clk          =>   b_mac_out[15]     ) = (0,0);
(clk          =>   b_mac_out[16]     ) = (0,0);
(clk          =>   b_mac_out[17]     ) = (0,0);
(clk          =>   b_mac_out[18]     ) = (0,0);
(clk          =>   b_mac_out[19]     ) = (0,0);
(clk          =>   b_mac_out[20]     ) = (0,0);
(clk          =>   b_mac_out[21]     ) = (0,0);
(clk          =>   b_mac_out[22]     ) = (0,0);
(clk          =>   b_mac_out[23]     ) = (0,0);
(clk          =>   a_overflow        ) = (0,0);
(a_dinx[0]    =>   a_mac_out[0]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[0]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[0]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[0]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[0]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[0]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[0]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[0]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[0]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[1]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[1]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[1]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[1]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[1]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[1]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[1]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[1]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[1]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[1]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[2]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[2]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[2]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[2]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[2]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[2]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[2]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[2]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[2]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[2]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[2]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[3]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[3]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[3]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[3]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[3]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[3]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[3]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[3]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[3]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[3]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[3]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[3]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[3]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[4]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[4]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[4]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[4]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[4]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[4]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[4]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[4]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[4]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[4]      ) = (0,0);
(b_dinx[4]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[4]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[4]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[4]      ) = (0,0);
(b_diny[1]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[4]      ) = (0,0);
(a_dinz[10]   =>   a_mac_out[4]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[4]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[5]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[5]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[5]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[5]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[5]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[5]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[5]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[5]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[5]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[5]      ) = (0,0);
(b_dinx[4]    =>   a_mac_out[5]      ) = (0,0);
(b_dinx[5]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[5]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[5]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[5]      ) = (0,0);
(b_diny[1]    =>   a_mac_out[5]      ) = (0,0);
(b_diny[2]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[5]      ) = (0,0);
(a_dinz[10]   =>   a_mac_out[5]      ) = (0,0);
(a_dinz[11]   =>   a_mac_out[5]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[5]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[6]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[4]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[5]    =>   a_mac_out[6]      ) = (0,0);
(b_dinx[6]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[6]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[6]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[6]      ) = (0,0);
(b_diny[1]    =>   a_mac_out[6]      ) = (0,0);
(b_diny[2]    =>   a_mac_out[6]      ) = (0,0);
(b_diny[3]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[6]      ) = (0,0);
(a_dinz[10]   =>   a_mac_out[6]      ) = (0,0);
(a_dinz[11]   =>   a_mac_out[6]      ) = (0,0);
(a_dinz[12]   =>   a_mac_out[6]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[6]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[6]    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[7]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[4]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[5]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[6]    =>   a_mac_out[7]      ) = (0,0);
(b_dinx[7]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[7]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[7]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[7]      ) = (0,0);
(b_diny[1]    =>   a_mac_out[7]      ) = (0,0);
(b_diny[2]    =>   a_mac_out[7]      ) = (0,0);
(b_diny[3]    =>   a_mac_out[7]      ) = (0,0);
(b_diny[4]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[7]      ) = (0,0);
(a_dinz[10]   =>   a_mac_out[7]      ) = (0,0);
(a_dinz[11]   =>   a_mac_out[7]      ) = (0,0);
(a_dinz[12]   =>   a_mac_out[7]      ) = (0,0);
(a_dinz[13]   =>   a_mac_out[7]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[7]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[6]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[7]    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[8]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[4]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[5]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[6]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[7]    =>   a_mac_out[8]      ) = (0,0);
(b_dinx[8]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[8]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[8]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[8]      ) = (0,0);
(b_diny[1]    =>   a_mac_out[8]      ) = (0,0);
(b_diny[2]    =>   a_mac_out[8]      ) = (0,0);
(b_diny[3]    =>   a_mac_out[8]      ) = (0,0);
(b_diny[4]    =>   a_mac_out[8]      ) = (0,0);
(b_diny[5]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[8]      ) = (0,0);
(a_dinz[10]   =>   a_mac_out[8]      ) = (0,0);
(a_dinz[11]   =>   a_mac_out[8]      ) = (0,0);
(a_dinz[12]   =>   a_mac_out[8]      ) = (0,0);
(a_dinz[13]   =>   a_mac_out[8]      ) = (0,0);
(a_dinz[14]   =>   a_mac_out[8]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[8]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[1]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[2]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[3]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[4]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[5]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[6]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[7]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[8]    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[9]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[0]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[1]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[2]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[3]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[4]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[5]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[6]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[7]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[8]    =>   a_mac_out[9]      ) = (0,0);
(b_dinx[9]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[0]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[1]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[2]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[3]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[4]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[5]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[6]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[7]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[8]    =>   a_mac_out[9]      ) = (0,0);
(a_diny[9]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[0]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[1]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[2]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[3]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[4]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[5]    =>   a_mac_out[9]      ) = (0,0);
(b_diny[6]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[0]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[1]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[2]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[3]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[4]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[5]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[6]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[7]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[8]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[9]    =>   a_mac_out[9]      ) = (0,0);
(a_dinz[10]   =>   a_mac_out[9]      ) = (0,0);
(a_dinz[11]   =>   a_mac_out[9]      ) = (0,0);
(a_dinz[12]   =>   a_mac_out[9]      ) = (0,0);
(a_dinz[13]   =>   a_mac_out[9]      ) = (0,0);
(a_dinz[14]   =>   a_mac_out[9]      ) = (0,0);
(a_dinz[15]   =>   a_mac_out[9]      ) = (0,0);
(a_dinz_en    =>   a_mac_out[9]      ) = (0,0);
(a_dinx[0]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[10]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[10]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[10]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[10]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[10]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[10]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[10]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[10]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[11]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[11]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[11]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[11]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[11]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[11]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[11]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[11]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[11]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[11]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[12]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[12]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[12]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[12]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[12]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[12]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[12]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[12]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[12]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[12]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[12]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[12]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[13]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[13]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[13]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[13]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[13]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[13]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[13]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[13]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[13]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[13]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[13]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[13]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[14]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[14]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[14]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[14]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[14]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[14]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[14]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[14]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[14]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[14]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[14]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[14]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[15]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[15]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[15]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[15]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[15]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[15]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[15]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[15]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[15]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[15]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[15]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[15]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[16]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[16]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[16]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[16]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[16]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[16]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[16]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[16]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[16]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[16]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[16]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[16]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[17]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[17]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[17]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[17]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[17]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[17]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[17]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[17]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[17]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[17]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[17]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[17]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[18]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[18]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[18]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[18]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[18]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[18]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[18]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[18]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[18]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[18]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[18]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[18]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[18]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[19]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[19]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[19]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[19]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[19]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[19]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[19]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[19]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[19]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[19]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[19]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[19]     ) = (0,0);
(b_dinz[1]    =>   a_mac_out[19]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[19]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[20]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[20]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[20]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[20]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[20]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[20]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[20]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[20]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[20]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[20]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[20]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[20]     ) = (0,0);
(b_dinz[1]    =>   a_mac_out[20]     ) = (0,0);
(b_dinz[2]    =>   a_mac_out[20]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[20]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[21]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[21]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[21]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[21]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[21]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[21]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[21]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[21]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[21]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[21]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[21]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[21]     ) = (0,0);
(b_dinz[1]    =>   a_mac_out[21]     ) = (0,0);
(b_dinz[2]    =>   a_mac_out[21]     ) = (0,0);
(b_dinz[3]    =>   a_mac_out[21]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[21]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[22]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[22]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[22]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[22]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[22]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[22]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[22]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[22]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[22]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[22]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[22]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[22]     ) = (0,0);
(b_dinz[1]    =>   a_mac_out[22]     ) = (0,0);
(b_dinz[2]    =>   a_mac_out[22]     ) = (0,0);
(b_dinz[3]    =>   a_mac_out[22]     ) = (0,0);
(b_dinz[4]    =>   a_mac_out[22]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[22]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[23]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[23]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[23]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[23]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[23]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[23]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[23]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[23]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[23]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[23]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[23]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[23]     ) = (0,0);
(b_dinz[1]    =>   a_mac_out[23]     ) = (0,0);
(b_dinz[2]    =>   a_mac_out[23]     ) = (0,0);
(b_dinz[3]    =>   a_mac_out[23]     ) = (0,0);
(b_dinz[4]    =>   a_mac_out[23]     ) = (0,0);
(b_dinz[5]    =>   a_mac_out[23]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[23]     ) = (0,0);
(a_dinx[0]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[1]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[2]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[3]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[4]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[5]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[6]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[7]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[8]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[9]    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[10]   =>   a_mac_out[24]     ) = (0,0);
(a_dinx[11]   =>   a_mac_out[24]     ) = (0,0);
(a_dinx[12]   =>   a_mac_out[24]     ) = (0,0);
(b_dinx[0]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[1]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[2]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[3]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[4]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[5]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[6]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[7]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[8]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[9]    =>   a_mac_out[24]     ) = (0,0);
(b_dinx[10]   =>   a_mac_out[24]     ) = (0,0);
(b_dinx[11]   =>   a_mac_out[24]     ) = (0,0);
(b_dinx[12]   =>   a_mac_out[24]     ) = (0,0);
(a_diny[0]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[1]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[2]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[3]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[4]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[5]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[6]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[7]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[8]    =>   a_mac_out[24]     ) = (0,0);
(a_diny[9]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[0]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[1]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[2]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[3]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[4]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[5]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[6]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[7]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[8]    =>   a_mac_out[24]     ) = (0,0);
(b_diny[9]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[0]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[1]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[2]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[3]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[4]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[5]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[6]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[7]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[8]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[9]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz[10]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[11]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[12]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[13]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[14]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[15]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[16]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[17]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[18]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[19]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[20]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[21]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[22]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[23]   =>   a_mac_out[24]     ) = (0,0);
(a_dinz[24]   =>   a_mac_out[24]     ) = (0,0);
(b_dinz[0]    =>   a_mac_out[24]     ) = (0,0);
(b_dinz[1]    =>   a_mac_out[24]     ) = (0,0);
(b_dinz[2]    =>   a_mac_out[24]     ) = (0,0);
(b_dinz[3]    =>   a_mac_out[24]     ) = (0,0);
(b_dinz[4]    =>   a_mac_out[24]     ) = (0,0);
(b_dinz[5]    =>   a_mac_out[24]     ) = (0,0);
(b_dinz[6]    =>   a_mac_out[24]     ) = (0,0);
(a_dinz_en    =>   a_mac_out[24]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[0]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[0]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[0]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[0]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[0]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[0]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[0]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[0]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[0]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[0]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[0]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[0]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[0]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[0]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[0]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[0]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[0]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[1]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[1]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[1]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[1]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[1]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[1]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[1]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[1]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[1]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[1]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[1]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[1]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[1]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[1]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[1]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[1]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[1]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[1]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[2]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[2]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[2]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[2]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[2]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[2]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[2]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[2]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[2]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[2]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[2]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[2]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[2]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[2]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[2]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[2]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[2]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[2]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[2]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[3]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[3]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[3]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[3]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[3]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[3]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[3]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[3]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[3]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[3]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[3]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[3]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[3]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[3]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[3]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[3]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[3]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[3]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[3]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[3]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[4]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[4]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[4]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[4]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[4]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[4]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[4]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[4]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[4]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[4]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[4]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[4]      ) = (0,0);
(b_dinz[7]    =>   b_mac_out[4]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[4]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[4]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[5]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[5]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[5]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[5]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[5]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[5]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[5]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[5]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[5]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[5]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[5]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[7]    =>   b_mac_out[5]      ) = (0,0);
(b_dinz[8]    =>   b_mac_out[5]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[5]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[5]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[6]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[6]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[6]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[6]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[6]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[6]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[6]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[6]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[6]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[6]      ) = (0,0);
(a_dinz[24]   =>   b_mac_out[6]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[7]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[8]    =>   b_mac_out[6]      ) = (0,0);
(b_dinz[9]    =>   b_mac_out[6]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[6]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[6]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[7]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[7]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[7]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[7]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[7]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[7]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[7]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[7]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[7]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[7]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz[24]   =>   b_mac_out[7]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[7]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[8]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[9]    =>   b_mac_out[7]      ) = (0,0);
(b_dinz[10]   =>   b_mac_out[7]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[7]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[7]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[8]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[8]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[8]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[8]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[8]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[8]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[8]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[8]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[8]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[8]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz[24]   =>   b_mac_out[8]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[7]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[8]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[9]    =>   b_mac_out[8]      ) = (0,0);
(b_dinz[10]   =>   b_mac_out[8]      ) = (0,0);
(b_dinz[11]   =>   b_mac_out[8]      ) = (0,0);
(b_dinz[21]   =>   b_mac_out[8]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[8]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[8]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[1]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[2]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[3]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[4]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[5]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[6]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[7]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[8]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[9]    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[10]   =>   b_mac_out[9]      ) = (0,0);
(a_dinx[11]   =>   b_mac_out[9]      ) = (0,0);
(a_dinx[12]   =>   b_mac_out[9]      ) = (0,0);
(b_dinx[0]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[1]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[2]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[3]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[4]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[5]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[6]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[7]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[8]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[9]    =>   b_mac_out[9]      ) = (0,0);
(b_dinx[10]   =>   b_mac_out[9]      ) = (0,0);
(b_dinx[11]   =>   b_mac_out[9]      ) = (0,0);
(b_dinx[12]   =>   b_mac_out[9]      ) = (0,0);
(a_diny[0]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[1]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[2]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[3]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[4]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[5]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[6]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[7]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[8]    =>   b_mac_out[9]      ) = (0,0);
(a_diny[9]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[0]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[1]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[2]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[3]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[4]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[5]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[6]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[7]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[8]    =>   b_mac_out[9]      ) = (0,0);
(b_diny[9]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[0]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[1]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[2]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[3]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[4]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[5]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[6]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[7]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[8]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[9]    =>   b_mac_out[9]      ) = (0,0);
(a_dinz[10]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[11]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[12]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[13]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[14]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[15]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[16]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[17]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[18]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[19]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[20]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[21]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[22]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[23]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz[24]   =>   b_mac_out[9]      ) = (0,0);
(b_dinz[0]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[1]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[2]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[3]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[4]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[5]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[6]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[7]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[8]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[9]    =>   b_mac_out[9]      ) = (0,0);
(b_dinz[10]   =>   b_mac_out[9]      ) = (0,0);
(b_dinz[11]   =>   b_mac_out[9]      ) = (0,0);
(b_dinz[12]   =>   b_mac_out[9]      ) = (0,0);
(a_dinz_en    =>   b_mac_out[9]      ) = (0,0);
(b_dinz_en    =>   b_mac_out[9]      ) = (0,0);
(a_dinx[0]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[10]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[10]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[10]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[10]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[10]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[10]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[10]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[10]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[10]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[10]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[10]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[10]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[10]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[10]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[10]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[10]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[10]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[10]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[11]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[11]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[11]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[11]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[11]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[11]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[11]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[11]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[11]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[11]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[11]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[11]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[11]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[11]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[11]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[11]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[11]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[11]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[11]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[12]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[12]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[12]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[12]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[12]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[12]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[12]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[12]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[12]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[12]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[12]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[12]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[12]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[12]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[12]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[12]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[12]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[12]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[12]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[12]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[13]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[13]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[13]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[13]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[13]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[13]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[13]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[13]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[13]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[13]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[13]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[13]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[13]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[13]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[13]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[14]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[14]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[14]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[14]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[14]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[14]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[14]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[14]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[14]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[14]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[14]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[14]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[14]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[14]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[14]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[15]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[15]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[15]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[15]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[15]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[15]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[15]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[15]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[15]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[15]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[15]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[15]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[15]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[15]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[15]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[16]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[16]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[16]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[16]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[16]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[16]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[16]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[16]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[16]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[16]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[16]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[16]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[16]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[16]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[16]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[17]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[17]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[17]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[17]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[17]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[17]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[17]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[17]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[17]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[17]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[17]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[17]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[17]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[17]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[17]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[18]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[18]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[18]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[18]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[18]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[18]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[18]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[18]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[18]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[18]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[18]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[18]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[18]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[18]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[18]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[19]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[19]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[19]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[19]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[19]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[19]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[19]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[19]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[19]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[19]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[19]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[19]     ) = (0,0);
(b_dinz[22]   =>   b_mac_out[19]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[19]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[19]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[20]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[20]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[20]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[20]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[20]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[20]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[20]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[20]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[20]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[20]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[20]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[22]   =>   b_mac_out[20]     ) = (0,0);
(b_dinz[23]   =>   b_mac_out[20]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[20]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[20]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[21]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[21]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[21]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[21]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[21]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[21]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[21]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[21]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[21]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[21]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[21]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[22]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[23]   =>   b_mac_out[21]     ) = (0,0);
(b_dinz[24]   =>   b_mac_out[21]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[21]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[21]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[22]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[22]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[22]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[22]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[22]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[22]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[22]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[22]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[22]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[22]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[22]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[22]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[23]   =>   b_mac_out[22]     ) = (0,0);
(b_dinz[24]   =>   b_mac_out[22]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[22]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[22]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[6]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[7]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[8]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[9]    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[10]   =>   b_mac_out[23]     ) = (0,0);
(a_dinx[11]   =>   b_mac_out[23]     ) = (0,0);
(a_dinx[12]   =>   b_mac_out[23]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[23]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[23]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[23]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[23]     ) = (0,0);
(a_diny[0]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[1]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[2]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[3]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[4]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[5]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[6]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[7]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[8]    =>   b_mac_out[23]     ) = (0,0);
(a_diny[9]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[23]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[0]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[1]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[2]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[3]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[4]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[5]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[6]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[7]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[8]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[9]    =>   b_mac_out[23]     ) = (0,0);
(a_dinz[10]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[11]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[12]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[13]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[14]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[15]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[16]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[17]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[18]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[19]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[20]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[21]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[22]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[23]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz[24]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[23]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[22]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[23]   =>   b_mac_out[23]     ) = (0,0);
(b_dinz[24]   =>   b_mac_out[23]     ) = (0,0);
(a_dinz_en    =>   b_mac_out[23]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[23]     ) = (0,0);
(a_dinx[0]    =>   b_mac_out[24]     ) = (0,0);
(a_dinx[1]    =>   b_mac_out[24]     ) = (0,0);
(a_dinx[2]    =>   b_mac_out[24]     ) = (0,0);
(a_dinx[3]    =>   b_mac_out[24]     ) = (0,0);
(a_dinx[4]    =>   b_mac_out[24]     ) = (0,0);
(a_dinx[5]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[0]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[1]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[2]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[3]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[4]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[5]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[6]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[7]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[8]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[9]    =>   b_mac_out[24]     ) = (0,0);
(b_dinx[10]   =>   b_mac_out[24]     ) = (0,0);
(b_dinx[11]   =>   b_mac_out[24]     ) = (0,0);
(b_dinx[12]   =>   b_mac_out[24]     ) = (0,0);
(b_diny[0]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[1]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[2]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[3]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[4]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[5]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[6]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[7]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[8]    =>   b_mac_out[24]     ) = (0,0);
(b_diny[9]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[0]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[1]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[2]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[3]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[4]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[5]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[6]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[7]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[8]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[9]    =>   b_mac_out[24]     ) = (0,0);
(b_dinz[10]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[11]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[12]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[13]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[14]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[15]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[16]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[17]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[18]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[19]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[20]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[21]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[22]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[23]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz[24]   =>   b_mac_out[24]     ) = (0,0);
(b_dinz_en    =>   b_mac_out[24]     ) = (0,0);
(a_dinx[0]    =>   a_overflow        ) = (0,0);
(a_dinx[1]    =>   a_overflow        ) = (0,0);
(a_dinx[2]    =>   a_overflow        ) = (0,0);
(a_dinx[3]    =>   a_overflow        ) = (0,0);
(a_dinx[4]    =>   a_overflow        ) = (0,0);
(a_dinx[5]    =>   a_overflow        ) = (0,0);
(a_dinx[6]    =>   a_overflow        ) = (0,0);
(a_dinx[7]    =>   a_overflow        ) = (0,0);
(a_dinx[8]    =>   a_overflow        ) = (0,0);
(a_dinx[9]    =>   a_overflow        ) = (0,0);
(a_dinx[10]   =>   a_overflow        ) = (0,0);
(a_dinx[11]   =>   a_overflow        ) = (0,0);
(a_dinx[12]   =>   a_overflow        ) = (0,0);
(b_dinx[0]    =>   a_overflow        ) = (0,0);
(b_dinx[1]    =>   a_overflow        ) = (0,0);
(b_dinx[2]    =>   a_overflow        ) = (0,0);
(b_dinx[3]    =>   a_overflow        ) = (0,0);
(b_dinx[4]    =>   a_overflow        ) = (0,0);
(b_dinx[5]    =>   a_overflow        ) = (0,0);
(b_dinx[6]    =>   a_overflow        ) = (0,0);
(b_dinx[7]    =>   a_overflow        ) = (0,0);
(b_dinx[8]    =>   a_overflow        ) = (0,0);
(b_dinx[9]    =>   a_overflow        ) = (0,0);
(b_dinx[10]   =>   a_overflow        ) = (0,0);
(b_dinx[11]   =>   a_overflow        ) = (0,0);
(b_dinx[12]   =>   a_overflow        ) = (0,0);
(a_diny[0]    =>   a_overflow        ) = (0,0);
(a_diny[1]    =>   a_overflow        ) = (0,0);
(a_diny[2]    =>   a_overflow        ) = (0,0);
(a_diny[3]    =>   a_overflow        ) = (0,0);
(a_diny[4]    =>   a_overflow        ) = (0,0);
(a_diny[5]    =>   a_overflow        ) = (0,0);
(a_diny[6]    =>   a_overflow        ) = (0,0);
(a_diny[7]    =>   a_overflow        ) = (0,0);
(a_diny[8]    =>   a_overflow        ) = (0,0);
(a_diny[9]    =>   a_overflow        ) = (0,0);
(b_diny[0]    =>   a_overflow        ) = (0,0);
(b_diny[1]    =>   a_overflow        ) = (0,0);
(b_diny[2]    =>   a_overflow        ) = (0,0);
(b_diny[3]    =>   a_overflow        ) = (0,0);
(b_diny[4]    =>   a_overflow        ) = (0,0);
(b_diny[5]    =>   a_overflow        ) = (0,0);
(b_diny[6]    =>   a_overflow        ) = (0,0);
(b_diny[7]    =>   a_overflow        ) = (0,0);
(b_diny[8]    =>   a_overflow        ) = (0,0);
(b_diny[9]    =>   a_overflow        ) = (0,0);
(a_dinz[0]    =>   a_overflow        ) = (0,0);
(a_dinz[1]    =>   a_overflow        ) = (0,0);
(a_dinz[2]    =>   a_overflow        ) = (0,0);
(a_dinz[3]    =>   a_overflow        ) = (0,0);
(a_dinz[4]    =>   a_overflow        ) = (0,0);
(a_dinz[5]    =>   a_overflow        ) = (0,0);
(a_dinz[6]    =>   a_overflow        ) = (0,0);
(a_dinz[7]    =>   a_overflow        ) = (0,0);
(a_dinz[8]    =>   a_overflow        ) = (0,0);
(a_dinz[9]    =>   a_overflow        ) = (0,0);
(a_dinz[10]   =>   a_overflow        ) = (0,0);
(a_dinz[11]   =>   a_overflow        ) = (0,0);
(a_dinz[12]   =>   a_overflow        ) = (0,0);
(a_dinz[13]   =>   a_overflow        ) = (0,0);
(a_dinz[14]   =>   a_overflow        ) = (0,0);
(a_dinz[15]   =>   a_overflow        ) = (0,0);
(a_dinz[16]   =>   a_overflow        ) = (0,0);
(a_dinz[17]   =>   a_overflow        ) = (0,0);
(a_dinz[18]   =>   a_overflow        ) = (0,0);
(a_dinz[19]   =>   a_overflow        ) = (0,0);
(a_dinz[20]   =>   a_overflow        ) = (0,0);
(a_dinz[21]   =>   a_overflow        ) = (0,0);
(a_dinz[22]   =>   a_overflow        ) = (0,0);
(a_dinz[23]   =>   a_overflow        ) = (0,0);
(a_dinz[24]   =>   a_overflow        ) = (0,0);
(b_dinz[0]    =>   a_overflow        ) = (0,0);
(b_dinz[1]    =>   a_overflow        ) = (0,0);
(b_dinz[2]    =>   a_overflow        ) = (0,0);
(b_dinz[3]    =>   a_overflow        ) = (0,0);
(b_dinz[4]    =>   a_overflow        ) = (0,0);
(b_dinz[5]    =>   a_overflow        ) = (0,0);
(b_dinz[6]    =>   a_overflow        ) = (0,0);
(b_dinz[7]    =>   a_overflow        ) = (0,0);
(b_dinz[8]    =>   a_overflow        ) = (0,0);
(b_dinz[9]    =>   a_overflow        ) = (0,0);
(b_dinz[10]   =>   a_overflow        ) = (0,0);
(b_dinz[11]   =>   a_overflow        ) = (0,0);
(b_dinz[12]   =>   a_overflow        ) = (0,0);
(b_dinz[13]   =>   a_overflow        ) = (0,0);
(b_dinz[14]   =>   a_overflow        ) = (0,0);
(b_dinz[15]   =>   a_overflow        ) = (0,0);
(b_dinz[16]   =>   a_overflow        ) = (0,0);
(b_dinz[17]   =>   a_overflow        ) = (0,0);
(b_dinz[18]   =>   a_overflow        ) = (0,0);
(b_dinz[19]   =>   a_overflow        ) = (0,0);
(b_dinz[20]   =>   a_overflow        ) = (0,0);
(b_dinz[21]   =>   a_overflow        ) = (0,0);
(b_dinz[22]   =>   a_overflow        ) = (0,0);
(b_dinz[23]   =>   a_overflow        ) = (0,0);
(a_dinz_en    =>   a_overflow        ) = (0,0);
(a_dinx[0]    =>   b_overflow        ) = (0,0);
(a_dinx[1]    =>   b_overflow        ) = (0,0);
(a_dinx[2]    =>   b_overflow        ) = (0,0);
(a_dinx[3]    =>   b_overflow        ) = (0,0);
(a_dinx[4]    =>   b_overflow        ) = (0,0);
(a_dinx[5]    =>   b_overflow        ) = (0,0);
(b_dinx[0]    =>   b_overflow        ) = (0,0);
(b_dinx[1]    =>   b_overflow        ) = (0,0);
(b_dinx[2]    =>   b_overflow        ) = (0,0);
(b_dinx[3]    =>   b_overflow        ) = (0,0);
(b_dinx[4]    =>   b_overflow        ) = (0,0);
(b_dinx[5]    =>   b_overflow        ) = (0,0);
(b_dinx[6]    =>   b_overflow        ) = (0,0);
(b_dinx[7]    =>   b_overflow        ) = (0,0);
(b_dinx[8]    =>   b_overflow        ) = (0,0);
(b_dinx[9]    =>   b_overflow        ) = (0,0);
(b_dinx[10]   =>   b_overflow        ) = (0,0);
(b_dinx[11]   =>   b_overflow        ) = (0,0);
(b_dinx[12]   =>   b_overflow        ) = (0,0);
(b_diny[0]    =>   b_overflow        ) = (0,0);
(b_diny[1]    =>   b_overflow        ) = (0,0);
(b_diny[2]    =>   b_overflow        ) = (0,0);
(b_diny[3]    =>   b_overflow        ) = (0,0);
(b_diny[4]    =>   b_overflow        ) = (0,0);
(b_diny[5]    =>   b_overflow        ) = (0,0);
(b_diny[6]    =>   b_overflow        ) = (0,0);
(b_diny[7]    =>   b_overflow        ) = (0,0);
(b_diny[8]    =>   b_overflow        ) = (0,0);
(b_diny[9]    =>   b_overflow        ) = (0,0);
(b_dinz[0]    =>   b_overflow        ) = (0,0);
(b_dinz[1]    =>   b_overflow        ) = (0,0);
(b_dinz[2]    =>   b_overflow        ) = (0,0);
(b_dinz[3]    =>   b_overflow        ) = (0,0);
(b_dinz[4]    =>   b_overflow        ) = (0,0);
(b_dinz[5]    =>   b_overflow        ) = (0,0);
(b_dinz[6]    =>   b_overflow        ) = (0,0);
(b_dinz[7]    =>   b_overflow        ) = (0,0);
(b_dinz[8]    =>   b_overflow        ) = (0,0);
(b_dinz[9]    =>   b_overflow        ) = (0,0);
(b_dinz[10]   =>   b_overflow        ) = (0,0);
(b_dinz[11]   =>   b_overflow        ) = (0,0);
(b_dinz[12]   =>   b_overflow        ) = (0,0);
(b_dinz[13]   =>   b_overflow        ) = (0,0);
(b_dinz[14]   =>   b_overflow        ) = (0,0);
(b_dinz[15]   =>   b_overflow        ) = (0,0);
(b_dinz[16]   =>   b_overflow        ) = (0,0);
(b_dinz[17]   =>   b_overflow        ) = (0,0);
(b_dinz[18]   =>   b_overflow        ) = (0,0);
(b_dinz[19]   =>   b_overflow        ) = (0,0);
(b_dinz[20]   =>   b_overflow        ) = (0,0);
(b_dinz[21]   =>   b_overflow        ) = (0,0);
(b_dinz[22]   =>   b_overflow        ) = (0,0);
(b_dinz[23]   =>   b_overflow        ) = (0,0);
(b_dinz[24]   =>   b_overflow        ) = (0,0);
(b_dinz_en    =>   b_overflow        ) = (0,0);


//timingcheck
$setuphold(posedge clk,    a_dinx[0] , 0,0); 
$setuphold(posedge clk,    a_dinx[1] , 0,0); 
$setuphold(posedge clk,    a_dinx[10], 0,0);  
$setuphold(posedge clk,    a_dinx[11], 0,0);  
$setuphold(posedge clk,    a_dinx[12], 0,0); 
$setuphold(posedge clk,    a_dinx[2] , 0,0); 
$setuphold(posedge clk,    a_dinx[3] , 0,0); 
$setuphold(posedge clk,    a_dinx[4] , 0,0);  
$setuphold(posedge clk,    a_dinx[5] , 0,0);  
$setuphold(posedge clk,    a_dinx[6] , 0,0);  
$setuphold(posedge clk,    a_dinx[7] , 0,0); 
$setuphold(posedge clk,    a_dinx[8] , 0,0); 
$setuphold(posedge clk,    a_dinx[9] , 0,0);  
$setuphold(posedge clk,    a_diny[0] , 0,0);  
$setuphold(posedge clk,    a_diny[1] , 0,0);  
$setuphold(posedge clk,    a_diny[2] , 0,0);  
$setuphold(posedge clk,    a_diny[3] , 0,0); 
$setuphold(posedge clk,    a_diny[4] , 0,0);  
$setuphold(posedge clk,    a_diny[5] , 0,0);  
$setuphold(posedge clk,    a_diny[6] , 0,0);  
$setuphold(posedge clk,    a_diny[7] , 0,0);  
$setuphold(posedge clk,    a_diny[8] , 0,0);  
$setuphold(posedge clk,    a_diny[9] , 0,0);  
$setuphold(posedge clk,    a_dinz[0] , 0,0); 
$setuphold(posedge clk,    a_dinz[1] , 0,0);  
$setuphold(posedge clk,    a_dinz[10], 0,0); 
$setuphold(posedge clk,    a_dinz[11], 0,0); 
$setuphold(posedge clk,    a_dinz[12], 0,0); 
$setuphold(posedge clk,    a_dinz[13], 0,0);  
$setuphold(posedge clk,    a_dinz[14], 0,0); 
$setuphold(posedge clk,    a_dinz[15], 0,0);  
$setuphold(posedge clk,    a_dinz[16], 0,0); 
$setuphold(posedge clk,    a_dinz[17], 0,0);  
$setuphold(posedge clk,    a_dinz[18], 0,0);  
$setuphold(posedge clk,    a_dinz[19], 0,0);   
$setuphold(posedge clk,    a_dinz[2] , 0,0);  
$setuphold(posedge clk,    a_dinz[20], 0,0);   
$setuphold(posedge clk,    a_dinz[21], 0,0); 
$setuphold(posedge clk,    a_dinz[22], 0,0); 
$setuphold(posedge clk,    a_dinz[23], 0,0); 
$setuphold(posedge clk,    a_dinz[24], 0,0); 
$setuphold(posedge clk,    a_dinz[3] , 0,0);  
$setuphold(posedge clk,    a_dinz[4] , 0,0);  
$setuphold(posedge clk,    a_dinz[5] , 0,0); 
$setuphold(posedge clk,    a_dinz[6] , 0,0); 
$setuphold(posedge clk,    a_dinz[7] , 0,0); 
$setuphold(posedge clk,    a_dinz[8] , 0,0); 
$setuphold(posedge clk,    a_dinz[9] , 0,0); 
$setuphold(posedge clk,    a_dinz_en , 0,0);  
$setuphold(posedge clk,    a_mac_out_cen ,0,0);
$setuphold(posedge clk,    a_out_sr   ,0,0);
$setuphold(posedge clk,    b_dinx[0]  ,0,0);  
$setuphold(posedge clk,    b_dinx[1]  ,0,0); 
$setuphold(posedge clk,    b_dinx[10] ,0,0);  
$setuphold(posedge clk,    b_dinx[11] ,0,0); 
$setuphold(posedge clk,    b_dinx[12] ,0,0); 
$setuphold(posedge clk,    b_dinx[2]  ,0,0); 
$setuphold(posedge clk,    b_dinx[3]  ,0,0); 
$setuphold(posedge clk,    b_dinx[4]  ,0,0); 
$setuphold(posedge clk,    b_dinx[5]  ,0,0); 
$setuphold(posedge clk,    b_dinx[6]  ,0,0); 
$setuphold(posedge clk,    b_dinx[7]  ,0,0); 
$setuphold(posedge clk,    b_dinx[8]  ,0,0); 
$setuphold(posedge clk,    b_dinx[9]  ,0,0); 
$setuphold(posedge clk,    b_diny[0]  ,0,0); 
$setuphold(posedge clk,    b_diny[1]  ,0,0); 
$setuphold(posedge clk,    b_diny[2]  ,0,0); 
$setuphold(posedge clk,    b_diny[3]  ,0,0); 
$setuphold(posedge clk,    b_diny[4]  ,0,0); 
$setuphold(posedge clk,    b_diny[5]  ,0,0); 
$setuphold(posedge clk,    b_diny[6]  ,0,0); 
$setuphold(posedge clk,    b_diny[7]  ,0,0); 
$setuphold(posedge clk,    b_diny[8]  ,0,0);  
$setuphold(posedge clk,    b_diny[9]  ,0,0); 
$setuphold(posedge clk,    b_dinz[0]  ,0,0); 
$setuphold(posedge clk,    b_dinz[1]  ,0,0); 
$setuphold(posedge clk,    b_dinz[10] ,0,0); 
$setuphold(posedge clk,    b_dinz[11] ,0,0); 
$setuphold(posedge clk,    b_dinz[12] ,0,0);  
$setuphold(posedge clk,    b_dinz[13] ,0,0); 
$setuphold(posedge clk,    b_dinz[14] ,0,0); 
$setuphold(posedge clk,    b_dinz[15] ,0,0); 
$setuphold(posedge clk,    b_dinz[16] ,0,0); 
$setuphold(posedge clk,    b_dinz[17] ,0,0); 
$setuphold(posedge clk,    b_dinz[18] ,0,0); 
$setuphold(posedge clk,    b_dinz[19] ,0,0); 
$setuphold(posedge clk,    b_dinz[2]  ,0,0);   
$setuphold(posedge clk,    b_dinz[20] ,0,0); 
$setuphold(posedge clk,    b_dinz[21] ,0,0); 
$setuphold(posedge clk,    b_dinz[22] ,0,0);  
$setuphold(posedge clk,    b_dinz[23] ,0,0);  
$setuphold(posedge clk,    b_dinz[3]  ,0,0); 
$setuphold(posedge clk,    b_dinz[4]  ,0,0); 
$setuphold(posedge clk,    b_dinz[5]  ,0,0); 
$setuphold(posedge clk,    b_dinz[6]  ,0,0); 
$setuphold(posedge clk,    b_dinz[7]  ,0,0); 
$setuphold(posedge clk,    b_dinz[8]  ,0,0); 
$setuphold(posedge clk,    b_dinz[9]  ,0,0); 
		endspecify

endmodule
module mac_dff_sync(q,clk,d,rstn,setn,cen);
input clk;
input d;
input rstn;
input setn;
input cen;
output q;
reg q;
always@(posedge clk)
begin
  if(!rstn)
    q <= 1'b0;
  else if(!setn)
    q <= 1'b1;
  else if(cen)
    q <= d;
end

endmodule

module mac_dff_async(q,clk,d,rstn,setn,cen);
input clk;
input d;
input rstn;   
input setn;   
input cen;    
output q;
reg q;
always@(posedge clk or negedge rstn or negedge setn)                                  
begin
  if(!rstn)   
    q <= 1'b0;
  else if(!setn)   
    q <= 1'b1;
  else if(cen)
    q <= d;   
end

endmodule

///////////// H6_BASIC_IO simulation model ///////////////

module H6_BASIC_IO(
     in
    ,f_oen
    ,f_out
    ,PAD
);

output       in;
input        f_oen;
input        f_out;
inout        PAD;

parameter    cfg_out_sel              = 2'b00;   // 00:1   01:0   10: out   11:~out
parameter    cfg_oen_sel              = 2'b00;   // 00:1   01:0   10: oen   11:~oen
parameter    cfg_keep                 = 2'b00; //pullup/pulldown/keep
parameter    cfg_ds                   = 1'b0;  //for drive strenth
parameter    cfg_nc                   = 1'b0;  //reserved

//reg PAD_reg;
wire out_en;
wire out_data;

assign in = PAD;
assign out_en = (cfg_oen_sel == 2'b00) ? 1'b1 :
				(cfg_oen_sel == 2'b01) ? 1'b0 :
				(cfg_oen_sel == 2'b10) ? f_oen :
				(cfg_oen_sel == 2'b11) ? ~f_oen : 1'bx; 
				
assign out_data = (cfg_out_sel == 2'b00) ? 1'b1 :
				  (cfg_out_sel == 2'b01) ? 1'b0 :
				  (cfg_out_sel == 2'b10) ? f_out :
				  (cfg_out_sel == 2'b11) ? ~f_out : 1'bx; 

				  
assign PAD = ~out_en ? out_data : 1'bz;
//always@(out_en or out_data)
//begin
//if(!out_en)
//    PAD_reg = out_data;
//else
//    PAD_reg= 1'bz;
//end
//
//assign PAD = PAD_reg; 
endmodule

///////////// H6_IOC_FUN simulation model ///////////////
module H6_IOC_FUN(
     clk_en
    ,oen
    ,f_oen
    ,out
    ,f_out
    ,f_out_fb
    ,in
    ,f_in
    ,ioc_clk_out
    ,clkfb
    ,fclk
    ,rstn
    ,setn
);

input          clk_en;
input          oen;
output         f_oen;
input  [1:0]   out;
output         f_out;
output         f_out_fb;
input          in;
output [1:0]   f_in;
output	       ioc_clk_out;
input          fclk;
input          clkfb;
input          rstn;
input          setn;

parameter cfg_nc             = 1'b0;
parameter cfg_ddr            = 1'b0;
parameter cfg_foen_sel       = 1'b0;
parameter cfg_fout_sel       = 1'b0;
parameter cfg_fin_sel        = 1'b0;
parameter cfg_fclk_inv       = 1'b0;
parameter cfg_fclk_gate_en   = 1'b0;
parameter cfg_setn_inv       = 1'b0;
parameter cfg_setn_sync      = 1'b0;
parameter cfg_oen_setn_en    = 1'b0;
parameter cfg_od_setn_en     = 1'b0;
parameter cfg_id_setn_en     = 1'b0;
parameter cfg_rstn_inv       = 1'b0;
parameter cfg_rstn_sync      = 1'b0;
parameter cfg_oen_rstn_en    = 1'b0;
parameter cfg_od_rstn_en     = 1'b0;
parameter cfg_id_rstn_en     = 1'b0;

//SIMULATION Model
`ifndef DLY
    `define DLY #1
`endif

reg cf_rstn;
initial begin
    cf_rstn = 1'b0;
    #1;
    cf_rstn = 1'b1;
end
//wire fclk_inv_cfg = cfg_fclk_inv ? ~fclk : fclk;
wire fclk_inv_cfg = fclk;
wire rstn_inv_cfg = cfg_rstn_inv ? ~rstn : rstn;
wire setn_inv_cfg = cfg_setn_inv ? ~setn : setn;

reg  fclk_gate_en = cfg_fclk_gate_en;
wire fclk_gate;
wire fclk_gate_mux;

ioc_dff_ar rstn_syn (
     .ck    (fclk_gate_mux )
    ,.d     (rstn_inv_cfg  )
    ,.q     (rstn_reg      )
    ,.rstn  (cf_rstn       )
);

ioc_dff_ar setn_syn (
     .ck    (fclk_gate_mux )
    ,.d     (setn_inv_cfg  )
    ,.q     (setn_reg      )
    ,.rstn  (cf_rstn       )
);

assign rstn_reg_mux = cfg_rstn_sync ? rstn_inv_cfg | rstn_reg : rstn_inv_cfg;
assign setn_reg_mux = cfg_setn_sync ? setn_inv_cfg | setn_reg : setn_inv_cfg;

assign oen_rstn = cfg_oen_rstn_en ? rstn_reg_mux : 1'b1;
assign od_rstn  = cfg_od_rstn_en ? rstn_reg_mux : 1'b1;
assign id_rstn  = cfg_id_rstn_en ? rstn_reg_mux : 1'b1;

assign t_oen_setn = cfg_oen_setn_en ? setn_reg_mux : 1'b1;
assign t_od_setn  = cfg_od_setn_en ? setn_reg_mux : 1'b1;
assign t_id_setn  = cfg_id_setn_en ? setn_reg_mux : 1'b1;

assign oen_setn = cf_rstn & t_oen_setn;
assign od_setn  = cf_rstn & t_od_setn;
assign id_setn  = cf_rstn & t_id_setn;

always@(*)
begin
    if (cfg_fclk_gate_en)
        fclk_gate_en <= 1'b1;
    else
    begin
        if (!fclk_inv_cfg)
            fclk_gate_en <= clk_en;
        else
            fclk_gate_en <= fclk_gate_en;
    end
end

assign fclk_gate_mux = fclk_gate_en & fclk_inv_cfg;
assign ioc_clk_out = clkfb;

ioc_dff_asr u0_oen(
     .ck     ( fclk_gate_mux )
    ,.d      ( oen           )
    ,.q      ( oen_reg       )
    ,.rstn   ( oen_rstn      )
    ,.setn   ( oen_setn      )
);

ioc_dff_asr u1_oen(
     .ck     (~fclk_gate_mux )
    ,.d      ( oen           )
    ,.q      ( oen_regn      )
    ,.rstn   ( oen_rstn      )
    ,.setn   ( oen_setn      )
);

assign f_oen_sel = cfg_nc ? oen_regn : oen_reg;
assign f_oen = !cfg_foen_sel ? f_oen_sel : oen;

ioc_dff_asr u_od0(
     .ck     ( fclk_gate_mux )
    ,.d      ( out[0]        )
    ,.q      ( out_reg0      )
    ,.rstn   ( od_rstn       )
    ,.setn   ( od_setn       )
);

ioc_dffn_asr u_od1(
     .ckb    ( fclk_gate_mux )
    ,.d      ( out[1]        )
    ,.q      ( out_reg1      )
    ,.rstn   ( od_rstn       )
    ,.setn   ( od_setn       )
);

//assign ddr_sel = ~(fclk_gate_mux & cfg_ddr);
assign ddr_sel = ~(~(fclk_gate_mux & cfg_ddr) & cfg_fclk_inv);
assign f_out_ddr = ddr_sel ? out_reg1 : out_reg0;
assign f_out = !cfg_fout_sel ? f_out_ddr : out[0];
assign f_out_fb = f_out;

ioc_dff_asr u_id0(
     .ck     ( fclk_gate_mux )
    ,.d      ( in            )
    ,.q      ( in_reg0       )
    ,.rstn   ( id_rstn       )
    ,.setn   ( id_setn       )
);

ioc_dffn_asr u_id1(
     .ckb    ( fclk_gate_mux )
    ,.d      ( in            )
    ,.q      ( in_reg1       )
    ,.rstn   ( id_rstn       )
    ,.setn   ( id_setn       )
);

assign f_in[0] = !cfg_fin_sel ? in_reg0 : in;
assign f_in[1] = in_reg1;

endmodule

module ioc_dff_ar(
     ck
    ,d
    ,q
    ,rstn
);

input  ck;
input  d;
output q;
input  rstn;

reg q;

always@(posedge ck or negedge rstn)
begin
    if(~rstn)
        q <= `DLY 1'b0;
    else
        q <= `DLY d;
end

endmodule

module IOC_LVDS_v2 (
	//port
	geclk0_up_il,
	geclk0_up_ol,
	rxd_dr,
	txd_out,
	ted_out,
	shiftout0_il,
	shiftout0_ol,
	shiftout1_il,
	shiftout1_ol,
	q,

	oen,
	rxd_in,
	shiftin0_il,
	shiftin0_ol,
	shiftin1_il,
	shiftin1_ol,
	update_il,
	update_b_il,
	update_ol,
	update_b_ol,
	clken,
	rstn,
	setn,
	feclk,
	sclk,
	test,
	d,
    in_del,
    out_del,
    in_del_update,
    out_del_update,
    idel_update_o,
    odel_update_o
	//PARAMETER
	`ifdef FM_HACK
	,CFG_CK_INV
	,CFG_CK_PAD_EN
	,CFG_DDR_IN_NREG
	,CFG_DDR_IN_NREG_DFF
	,CFG_DDR_IN_PREG
	,CFG_DDR_IN_PREG_DFF
	,CFG_DDR_OUT
	,CFG_DDR_OUT_REG
	,CFG_DQS_CLK
	,CFG_ECLK_INV
	,CFG_FASTIN
	,CFG_FCLK_OUT_EN
	,CFG_FCLK0_I_EN
	,CFG_FCLK0_OEN
	,CFG_FCLK0_O_EN
	,CFG_FCLK0_RS_EN
	,CFG_FCLK0_UPI_EN
	,CFG_FCLK0_UPO_EN
	,CFG_FCLK1_I_EN
	,CFG_FCLK1_O_EN
	,CFG_FCLK_INV
	,CFG_FOUT_SEL
	,CFG_GEAR_IN
	,CFG_GEAR_OUT
	,CFG_GECLK0_I_EN
	,CFG_GECLK0_O_EN
	,CFG_GECLK1_I_EN
	,CFG_GECLK1_O_EN
	,CFG_GSCLK0_I_EN
	,CFG_GSCLK0_O_EN
	,CFG_GSCLK1_I_EN
	,CFG_GSCLK1_O_EN
	,CFG_IN_EN
	,CFG_OEN_INV
	,CFG_OEN_SEL
	,CFG_OFDBK
	,CFG_OUT_SEL
	,CFG_RSTN
	,CFG_SCLK_INV
	,CFG_SETN
	,CFG_SLAVE_IN
	,CFG_TEST
	`endif
	);
output	geclk0_up_il;
output	geclk0_up_ol;
output	rxd_dr;
output	txd_out;
output	ted_out;
output	shiftout0_il;
output	shiftout0_ol;
output	shiftout1_il;
output	shiftout1_ol;
output	[7:0]	q;

input	oen;
input	rxd_in;
input	shiftin0_il;
input	shiftin0_ol;
input	shiftin1_il;
input	shiftin1_ol;
input	update_il;
input	update_b_il;
input	update_ol;
input	update_b_ol;
input	clken;
input	rstn;
input	setn;
input	feclk;
input	sclk;
input	[7:0]	test;
input	[7:0]	d;

input [5:0]    in_del;
input [5:0]    out_del;
input    in_del_update;
input    out_del_update;
output [5:0]    idel_update_o;
output [5:0]    odel_update_o;

`ifdef FM_HACK
input	CFG_CK_INV;
input	CFG_CK_PAD_EN;
input	CFG_DDR_IN_NREG;
input	CFG_DDR_IN_NREG_DFF;
input	CFG_DDR_IN_PREG;
input	CFG_DDR_IN_PREG_DFF;
input	CFG_DDR_OUT;
input	CFG_DDR_OUT_REG;
input	CFG_DQS_CLK;
input	CFG_ECLK_INV;
input	CFG_FASTIN;
input	CFG_FCLK_OUT_EN;
input	CFG_FCLK0_I_EN;
input	CFG_FCLK0_OEN;
input	CFG_FCLK0_O_EN;
input	CFG_FCLK0_RS_EN;
input	CFG_FCLK0_UPI_EN;
input	CFG_FCLK0_UPO_EN;
input	CFG_FCLK1_I_EN;
input	CFG_FCLK1_O_EN;
input	CFG_FCLK_INV;
input	CFG_FOUT_SEL;
input	CFG_GEAR_OUT;
input	CFG_GECLK0_I_EN;
input	CFG_GECLK0_O_EN;
input	CFG_GECLK1_I_EN;
input	CFG_GECLK1_O_EN;
input	CFG_GSCLK0_I_EN;
input	CFG_GSCLK0_O_EN;
input	CFG_GSCLK1_I_EN;
input	CFG_GSCLK1_O_EN;
input	CFG_OEN_INV;
input	CFG_OFDBK;
input	CFG_SCLK_INV;
input	CFG_SLAVE_IN;
input	[7:0]	CFG_GEAR_IN;
input	[1:0]	CFG_IN_EN;
input	[3:0]	CFG_OEN_SEL;
input	[2:0]	CFG_OUT_SEL;
input	[4:0]	CFG_RSTN;
input	[4:0]	CFG_SETN;
input	[7:0]	CFG_TEST;
`else
parameter	CFG_CK_INV=1'b0;
parameter	CFG_CK_PAD_EN=1'b0;
parameter	CFG_DDR_IN_NREG=1'b0;
parameter	CFG_DDR_IN_NREG_DFF=1'b0;
parameter	CFG_DDR_IN_PREG=1'b0;
parameter	CFG_DDR_IN_PREG_DFF=1'b0;
parameter	CFG_DDR_OUT=1'b0;
parameter	CFG_DDR_OUT_REG=1'b0;
parameter	CFG_DQS_CLK=1'b0;
parameter	CFG_ECLK_INV=1'b0;
parameter	CFG_FASTIN=1'b0;
parameter	CFG_FCLK_OUT_EN=1'b0;
parameter	CFG_FCLK0_I_EN=1'b0;
parameter	CFG_FCLK0_OEN=1'b0;
parameter	CFG_FCLK0_O_EN=1'b0;
parameter	CFG_FCLK0_RS_EN=1'b0;
parameter	CFG_FCLK0_UPI_EN=1'b0;
parameter	CFG_FCLK0_UPO_EN=1'b0;
parameter	CFG_FCLK1_I_EN=1'b0;
parameter	CFG_FCLK1_O_EN=1'b0;
parameter	CFG_FCLK_INV=1'b0;
parameter	CFG_FOUT_SEL=1'b0;
parameter	CFG_GEAR_OUT=1'b0;
parameter	CFG_GECLK0_I_EN=1'b0;
parameter	CFG_GECLK0_O_EN=1'b0;
parameter	CFG_GECLK1_I_EN=1'b0;
parameter	CFG_GECLK1_O_EN=1'b0;
parameter	CFG_GSCLK0_I_EN=1'b0;
parameter	CFG_GSCLK0_O_EN=1'b0;
parameter	CFG_GSCLK1_I_EN=1'b0;
parameter	CFG_GSCLK1_O_EN=1'b0;
parameter	CFG_OEN_INV=1'b0;
parameter	CFG_OFDBK=1'b0;
parameter	CFG_SCLK_INV=1'b0;
parameter	CFG_SLAVE_IN=1'b0;
parameter	CFG_GEAR_IN=8'b0;
parameter	CFG_IN_EN=2'b0;
parameter	CFG_OEN_SEL=4'b0;
parameter	CFG_OUT_SEL=3'b0;
parameter	CFG_RSTN=5'b0;
parameter	CFG_SETN=5'b0;
parameter	CFG_TEST=8'b0;
`endif
wire	[7:0]	CFG_GEAR_IN_              = ~CFG_GEAR_IN;
wire	[1:0]	CFG_IN_EN_                = ~CFG_IN_EN;
wire	[2:0]	CFG_OUT_SEL_              = ~CFG_OUT_SEL;
wire	[4:0]	CFG_RSTN_                 = ~CFG_RSTN;
wire	[4:0]	CFG_SETN_                 = ~CFG_SETN;
wire	[7:0]	CFG_TEST_                 = ~CFG_TEST;
wire			CFG_CK_INV_               = ~CFG_CK_INV;
wire			CFG_DDR_IN_NREG_          = ~CFG_DDR_IN_NREG;
wire			CFG_DDR_IN_NREG_DFF_      = ~CFG_DDR_IN_NREG_DFF;
wire			CFG_DDR_IN_PREG_          = ~CFG_DDR_IN_PREG;
wire			CFG_DDR_IN_PREG_DFF_      = ~CFG_DDR_IN_PREG_DFF;
wire			CFG_DDR_OUT_REG_          = ~CFG_DDR_OUT_REG;
wire			CFG_DQS_CLK_              = ~CFG_DQS_CLK;
wire			CFG_FASTIN_               = ~CFG_FASTIN;
wire			CFG_FOUT_SEL_             = ~CFG_FOUT_SEL;
wire			CFG_GEAR_OUT_             = ~CFG_GEAR_OUT;
wire			CFG_OEN_INV_              = ~CFG_OEN_INV;
wire			CFG_OFDBK_                = ~CFG_OFDBK;
wire			CFG_SLAVE_IN_             = ~CFG_SLAVE_IN;
`ifndef FM_HACK
reg gbl_clear_b;

wire GSR;
glbsr glbsr_inst(.GSR(GSR));
initial begin
gbl_clear_b = 1'b0;
@(posedge GSR);
gbl_clear_b = 1'b1;
end
`else
wire gbl_clear_b = 1'b1;
`endif

assign rxd_dr = CFG_CK_PAD_EN & rxd_in;
wire	txd_in,txd_in_b;
wire	fclk0_ol;
assign txd_in_b = (CFG_FCLK_OUT_EN == 1'b1) ? ~fclk0_ol : ~txd_in;
assign txd_out =	({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b001_110) ? 1'b0 :
					({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b010_101) ? txd_in_b :
					({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b100_011) ? !txd_in_b :
					({CFG_OUT_SEL,CFG_OUT_SEL_} == 6'b000_111) ? 1'b1 : 1'bx;
wire	datain;
assign datain =	({CFG_OFDBK,CFG_OFDBK_} == 2'b01) ? rxd_in :
				({CFG_OFDBK,CFG_OFDBK_} == 2'b10) ? txd_in : 1'bx;
// VPERL: GENERATED_BEG


CLK_v1 Iclk (
	.CFG_CKEN_INV		(CFG_CK_INV),
	.CFG_CKEN_INV_		(CFG_CK_INV_),
	.CFG_FCLK0_I_EN		(CFG_FCLK0_I_EN),
	.CFG_FCLK0_OEN		(CFG_FCLK0_OEN),
	.CFG_FCLK0_O_EN		(CFG_FCLK0_O_EN),
	.CFG_FCLK0_RS_EN	(CFG_FCLK0_RS_EN),
	.CFG_FCLK0_UPI_EN	(CFG_FCLK0_UPI_EN),
	.CFG_FCLK0_UPO_EN	(CFG_FCLK0_UPO_EN),
	.CFG_FCLK1_I_EN		(CFG_FCLK1_I_EN),
	.CFG_FCLK1_O_EN		(CFG_FCLK1_O_EN),
	.CFG_GECLK0_I_EN	(CFG_GECLK0_I_EN),
	.CFG_GECLK0_O_EN	(CFG_GECLK0_O_EN),
	.CFG_GECLK1_I_EN	(CFG_GECLK1_I_EN),
	.CFG_GECLK1_O_EN	(CFG_GECLK1_O_EN),
	.CFG_GSCLK0_I_EN	(CFG_GSCLK0_I_EN),
	.CFG_GSCLK0_O_EN	(CFG_GSCLK0_O_EN),
	.CFG_GSCLK1_I_EN	(CFG_GSCLK1_I_EN),
	.CFG_GSCLK1_O_EN	(CFG_GSCLK1_O_EN),
	.CFG_RSTN_ID_EN		(CFG_RSTN[4]),
	.CFG_RSTN_ID_EN_	(CFG_RSTN_[4]),
	.CFG_RSTN_INV		(CFG_RSTN[1]),
	.CFG_RSTN_INV_		(CFG_RSTN_[1]),
	.CFG_RSTN_OD_EN		(CFG_RSTN[3]),
	.CFG_RSTN_OD_EN_	(CFG_RSTN_[3]),
	.CFG_RSTN_OEN_EN	(CFG_RSTN[2]),
	.CFG_RSTN_OEN_EN_	(CFG_RSTN_[2]),
	.CFG_RSTN_SYNC		(CFG_RSTN[0]),
	.CFG_RSTN_SYNC_		(CFG_RSTN_[0]),
	.CFG_SETN_ID_EN		(CFG_SETN[4]),
	.CFG_SETN_ID_EN_	(CFG_SETN_[4]),
	.CFG_SETN_INV		(CFG_SETN[1]),
	.CFG_SETN_INV_		(CFG_SETN_[1]),
	.CFG_SETN_OD_EN		(CFG_SETN[3]),
	.CFG_SETN_OD_EN_	(CFG_SETN_[3]),
	.CFG_SETN_OEN_EN	(CFG_SETN[2]),
	.CFG_SETN_OEN_EN_	(CFG_SETN_[2]),
	.CFG_SETN_SYNC		(CFG_SETN[0]),
	.CFG_SETN_SYNC_		(CFG_SETN_[0]),
	.CFG_SCLK_INV  		(CFG_SCLK_INV),
	.CFG_ECLK_INV  		(CFG_ECLK_INV),
	.setn			(setn),
	.rstn			(rstn),
	.clk_en			(clken),
	.sclk			(sclk),
	.feclk			(feclk),

	.fclk0_il		(fclk0_il),
	.fclk0_oen		(oen_fclk0),
	.fclk0_ol		(fclk0_ol),
	.fclk1_il		(fclk1_il),
	.fclk1_ol		(fclk1_ol),
	.geclk0_il		(geclk0_il),
	.geclk0_ol		(geclk0_ol),
	.geclk0_up_il		(geclk0_up_il),
	.geclk0_up_ol		(geclk0_up_ol),
	.geclk1_il		(geclk1_il),
	.geclk1_ol		(geclk1_ol),
	.gsclk0_il		(gsclk0_il),
	.gsclk0_ol		(gsclk0_ol),
	.gsclk1_il		(gsclk1_il),
	.gsclk1_ol		(gsclk1_ol),
	.id_rst			(id_rst),
	.id_setn		(id_set_),
	.od_rst			(od_rst),
	.od_setn		(od_set_),
	.oen_rst		(oen_rst),
	.oen_setn		(oen_set_) 
);

ILOGIC Iilg (
	.datain			(datain),
	.fclk0			(fclk0_il),
	.fclk1			(fclk1_il),
	.geclk0			(geclk0_il),
	.geclk1			(geclk1_il),
	.gsclk0			(gsclk0_il),
	.gsclk1			(gsclk1_il),
	.init_b			(1'b1),
	.rst			(id_rst),
	.set_			(id_set_),
	.shiftin0		(shiftin0_il),
	.shiftin1		(shiftin1_il),
	.update			(update_il),
	.update_		(update_b_il),
	.usermode		(gbl_clear_b),
	.test			(test[7:0]),
	.CFG_DDR_IN_NREG	(CFG_DDR_IN_NREG),
	.CFG_DDR_IN_NREG_DFF	(CFG_DDR_IN_NREG_DFF),
	.CFG_DDR_IN_PREG	(CFG_DDR_IN_PREG),
	.CFG_DDR_IN_PREG_DFF	(CFG_DDR_IN_PREG_DFF),
	.CFG_DQS_CLK		(CFG_DQS_CLK),
	.CFG_FASTIN		(CFG_FASTIN),
	.CFG_SLAVE_IN		(CFG_SLAVE_IN),
	.CFG_TEST		(CFG_TEST[7:0]),
	.CFG_IN_EN		(CFG_IN_EN[1:0]),
	.CFG_GEAR_IN		(CFG_GEAR_IN[7:0]),
	.CFG_DDR_IN_NREG_	(CFG_DDR_IN_NREG_),
	.CFG_DDR_IN_NREG_DFF_	(CFG_DDR_IN_NREG_DFF_),
	.CFG_DDR_IN_PREG_	(CFG_DDR_IN_PREG_),
	.CFG_DDR_IN_PREG_DFF_	(CFG_DDR_IN_PREG_DFF_),
	.CFG_DQS_CLK_		(CFG_DQS_CLK_),
	.CFG_FASTIN_		(CFG_FASTIN_),
	.CFG_SLAVE_IN_		(CFG_SLAVE_IN_),
	.CFG_TEST_		(CFG_TEST_[7:0]),
	.CFG_IN_EN_		(CFG_IN_EN_[1:0]),
	.CFG_GEAR_IN_		(CFG_GEAR_IN_[7:0]),

	.shiftout0		(shiftout0_il),
	.shiftout1		(shiftout1_il),
	.dataout		(q[7:0]) 
);

OLOGIC Iolg (
	.fclk0			(fclk0_ol),
	.fclk1			(fclk1_ol),
	.geclk0			(geclk0_ol),
	.geclk1			(geclk1_ol),
	.gsclk0			(gsclk0_ol),
	.gsclk1			(gsclk1_ol),
	.rst			(od_rst),
	.set_			(od_set_),
	.shiftin0		(shiftin0_ol),
	.shiftin1		(shiftin1_ol),
	.update			(update_ol),
	.update_		(update_b_ol),
	.usermode		(gbl_clear_b),
	.datain			(d[7:0]),
	.CFG_DDR_OUT		(CFG_DDR_OUT),
	.CFG_DDR_OUT_REG	(CFG_DDR_OUT_REG),
	.CFG_DDR_OUT_REG_	(CFG_DDR_OUT_REG_),
	.CFG_FCLK_INV		(CFG_FCLK_INV),
	.CFG_FOUT_SEL		(CFG_FOUT_SEL),
	.CFG_FOUT_SEL_		(CFG_FOUT_SEL_),
	.CFG_GEAR_OUT		(CFG_GEAR_OUT),
	.CFG_GEAR_OUT_		(CFG_GEAR_OUT_),

	.dataout		(txd_in),
	.shiftout0		(shiftout0_ol),
	.shiftout1		(shiftout1_ol) 
);

OENC_v1 Ioen (
	.clk		(oen_fclk0),
	.gbl_clear_b	(gbl_clear_b),
	.init_b		(1'b1),
	.oen		(oen),
	.rst		(oen_rst),
	.set_		(oen_set_),
	.CFG_OEN_INV	(CFG_OEN_INV),
	.CFG_OEN_INV_	(CFG_OEN_INV_),
	.CFG_OEN_SEL	(CFG_OEN_SEL[3:0]),

	.f_oen		(ted_out) 
);
// VPERL: GENERATED_END
endmodule

module CLK_v1 (
	fclk0_il,
	fclk0_oen,
	fclk0_ol,
	fclk1_il,
	fclk1_ol,
	geclk0_il,
	geclk0_ol,
	geclk0_up_il,
	geclk0_up_ol,
	geclk1_il,
	geclk1_ol,
	gsclk0_il,
	gsclk0_ol,
	gsclk1_il,
	gsclk1_ol,
	id_rst,
	id_setn,
	od_rst,
	od_setn,
	oen_rst,
	oen_setn,
	//PARAMETER 
	CFG_CKEN_INV,
	CFG_CKEN_INV_,
	CFG_FCLK0_I_EN,
	CFG_FCLK0_OEN,
	CFG_FCLK0_O_EN,
	CFG_FCLK0_RS_EN,
	CFG_FCLK0_UPI_EN,
	CFG_FCLK0_UPO_EN,
	CFG_FCLK1_I_EN,
	CFG_FCLK1_O_EN,
	CFG_GECLK0_I_EN,
	CFG_GECLK0_O_EN,
	CFG_GECLK1_I_EN,
	CFG_GECLK1_O_EN,
	CFG_GSCLK0_I_EN,
	CFG_GSCLK0_O_EN,
	CFG_GSCLK1_I_EN,
	CFG_GSCLK1_O_EN,
	CFG_RSTN_ID_EN,
	CFG_RSTN_ID_EN_,
	CFG_RSTN_INV,
	CFG_RSTN_INV_,
	CFG_RSTN_OD_EN,
	CFG_RSTN_OD_EN_,
	CFG_RSTN_OEN_EN,
	CFG_RSTN_OEN_EN_,
	CFG_RSTN_SYNC,
	CFG_RSTN_SYNC_,
	CFG_SETN_ID_EN,
	CFG_SETN_ID_EN_,
	CFG_SETN_INV,
	CFG_SETN_INV_,
	CFG_SETN_OD_EN,
	CFG_SETN_OD_EN_,
	CFG_SETN_OEN_EN,
	CFG_SETN_OEN_EN_,
	CFG_SETN_SYNC,
	CFG_SETN_SYNC_,
	CFG_SCLK_INV,
	CFG_ECLK_INV,
	//PARAMETER END
	setn,
	rstn,
	clk_en,
	sclk,
	feclk
	);
output	fclk0_il;
output	fclk0_oen;
output	fclk0_ol;
output	fclk1_il;
output	fclk1_ol;
output	geclk0_il;
output	geclk0_ol;
output	geclk0_up_il;
output	geclk0_up_ol;
output	geclk1_il;
output	geclk1_ol;
output	gsclk0_il;
output	gsclk0_ol;
output	gsclk1_il;
output	gsclk1_ol;
output	id_rst;
output	id_setn;
output	od_rst;
output	od_setn;
output	oen_rst;
output	oen_setn;
input	CFG_CKEN_INV;
input	CFG_CKEN_INV_;
input	CFG_FCLK0_I_EN;
input	CFG_FCLK0_OEN;
input	CFG_FCLK0_O_EN;
input	CFG_FCLK0_RS_EN;
input	CFG_FCLK0_UPI_EN;
input	CFG_FCLK0_UPO_EN;
input	CFG_FCLK1_I_EN;
input	CFG_FCLK1_O_EN;
input	CFG_GECLK0_I_EN;
input	CFG_GECLK0_O_EN;
input	CFG_GECLK1_I_EN;
input	CFG_GECLK1_O_EN;
input	CFG_GSCLK0_I_EN;
input	CFG_GSCLK0_O_EN;
input	CFG_GSCLK1_I_EN;
input	CFG_GSCLK1_O_EN;
input	CFG_RSTN_ID_EN;
input	CFG_RSTN_ID_EN_;
input	CFG_RSTN_INV;
input	CFG_RSTN_INV_;
input	CFG_RSTN_OD_EN;
input	CFG_RSTN_OD_EN_;
input	CFG_RSTN_OEN_EN;
input	CFG_RSTN_OEN_EN_;
input	CFG_RSTN_SYNC;
input	CFG_RSTN_SYNC_;
input	CFG_SETN_ID_EN;
input	CFG_SETN_ID_EN_;
input	CFG_SETN_INV;
input	CFG_SETN_INV_;
input	CFG_SETN_OD_EN;
input	CFG_SETN_OD_EN_;
input	CFG_SETN_OEN_EN;
input	CFG_SETN_OEN_EN_;
input	CFG_SETN_SYNC;
input	CFG_SETN_SYNC_;
input	CFG_SCLK_INV;
input	CFG_ECLK_INV;
input	setn;
input	rstn;
input	clk_en;
input	sclk;
input	feclk;

wire ck_inv = ({CFG_CKEN_INV,CFG_CKEN_INV_} == 2'b01) ? clk_en :
			  ({CFG_CKEN_INV,CFG_CKEN_INV_} == 2'b10) ? ~clk_en : 1'b0;
wire sckinv = CFG_SCLK_INV ? ~sclk  : sclk;
wire eckinv = CFG_ECLK_INV ? ~feclk : feclk;
wire sclk_b,eclk_b;
reg	sck_reg,eck_reg;
always @(sckinv or ck_inv)
	if(sckinv == 0) sck_reg <= ck_inv;
always @(eckinv or ck_inv)
	if(eckinv == 0) eck_reg <= ck_inv;
assign sclk_b = (sckinv & sck_reg);
assign eclk_b = (eckinv & eck_reg);

wire fclk0_sr;
assign fclk0_sr = CFG_FCLK0_RS_EN & eclk_b;
assign geclk0_up_il = CFG_FCLK0_UPI_EN & eclk_b;
assign geclk0_up_ol = CFG_FCLK0_UPO_EN & eclk_b;
assign fclk0_oen = CFG_FCLK0_OEN & eclk_b;
assign geclk0_il = CFG_GECLK0_I_EN & eclk_b;
assign geclk1_il = CFG_GECLK1_I_EN & eclk_b;
assign fclk0_il = CFG_FCLK0_I_EN & eclk_b;
assign fclk1_il = CFG_FCLK1_I_EN & eclk_b;
assign geclk0_ol = CFG_GECLK0_O_EN & eclk_b;
assign geclk1_ol = CFG_GECLK1_O_EN & eclk_b;
assign fclk0_ol = CFG_FCLK0_O_EN & eclk_b;
assign fclk1_ol = CFG_FCLK1_O_EN & eclk_b;
assign gsclk0_ol = CFG_GSCLK0_O_EN & sclk_b;
assign gsclk1_ol = CFG_GSCLK1_O_EN & sclk_b;
assign gsclk0_il = CFG_GSCLK0_I_EN & sclk_b;
assign gsclk1_il = CFG_GSCLK1_I_EN & sclk_b;

wire set_inv = ({CFG_SETN_INV,CFG_SETN_INV_} == 2'b01) ? ~setn :
			   ({CFG_SETN_INV,CFG_SETN_INV_} == 2'b10) ? setn : 1'b0;
reg	set_reg;
always @(set_inv or fclk0_sr)
	if(fclk0_sr == 0) set_reg <= set_inv;
wire set_sync = (set_reg & fclk0_sr);
wire set_sel = ({CFG_SETN_SYNC,CFG_SETN_SYNC_} == 2'b01) ? set_inv :
			   ({CFG_SETN_SYNC,CFG_SETN_SYNC_} == 2'b10) ? set_sync : 1'b0;
wire od_set = ({CFG_SETN_OD_EN,CFG_SETN_OD_EN_} == 2'b01) ? 1'b1 :
			  ({CFG_SETN_OD_EN,CFG_SETN_OD_EN_} == 2'b10) ? ~set_sel : 1'b0;
wire id_set = ({CFG_SETN_ID_EN,CFG_SETN_ID_EN_} == 2'b01) ? 1'b1 :
			  ({CFG_SETN_ID_EN,CFG_SETN_ID_EN_} == 2'b10) ? ~set_sel : 1'b0;
wire oen_set = ({CFG_SETN_OEN_EN,CFG_SETN_OEN_EN_} == 2'b01) ? 1'b1 :
			   ({CFG_SETN_OEN_EN,CFG_SETN_OEN_EN_} == 2'b10) ? ~set_sel : 1'b0;
assign od_setn = od_set;
assign id_setn = id_set;
assign oen_setn = oen_set;
wire rst_inv = ({CFG_RSTN_INV,CFG_RSTN_INV_} == 2'b01) ? ~rstn :
			   ({CFG_RSTN_INV,CFG_RSTN_INV_} == 2'b10) ? rstn : 1'b0;
reg	rst_reg;
always @(rst_inv or fclk0_sr)
	if(fclk0_sr == 0) rst_reg <= rst_inv;
wire rst_sync = (rst_reg & fclk0_sr);
wire rst_sel = ({CFG_RSTN_SYNC,CFG_RSTN_SYNC_} == 2'b01) ? rst_inv :
			   ({CFG_RSTN_SYNC,CFG_RSTN_SYNC_} == 2'b10) ? rst_sync : 1'b0;
wire od_rst = ({CFG_RSTN_OD_EN,CFG_RSTN_OD_EN_} == 2'b01) ? 1'b0 :
			  ({CFG_RSTN_OD_EN,CFG_RSTN_OD_EN_} == 2'b10) ? rst_sel : 1'b1;
wire id_rst = ({CFG_RSTN_ID_EN,CFG_RSTN_ID_EN_} == 2'b01) ? 1'b0 :
			  ({CFG_RSTN_ID_EN,CFG_RSTN_ID_EN_} == 2'b10) ? rst_sel : 1'b1;
wire oen_rst = ({CFG_RSTN_OEN_EN,CFG_RSTN_OEN_EN_} == 2'b01) ? 1'b0 :
			   ({CFG_RSTN_OEN_EN,CFG_RSTN_OEN_EN_} == 2'b10) ? rst_sel : 1'b1;

endmodule

module OENC_v1 (
	f_oen,
	clk,
	gbl_clear_b,
	init_b,
	oen,
	rst,
	set_,
	CFG_OEN_INV,
	CFG_OEN_INV_,
	CFG_OEN_SEL
	);
output	f_oen;
input	clk,gbl_clear_b,init_b,oen,rst,set_;
input	CFG_OEN_INV;
input	CFG_OEN_INV_;
input	[3:0]	CFG_OEN_SEL;

wire	oen_inv;
assign oen_inv =({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b011) ? ~oen : 
				({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b101) ? oen :
				({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b000) ? 1'b0 :
				({CFG_OEN_INV,CFG_OEN_INV_,init_b} == 3'b001) ? 1'b0 : 1'bx;
reg		oen_psync;
reg		oen_nsync;

always @(posedge clk or posedge rst or negedge set_)
	if(~set_) oen_psync <= 1;
	else if(rst) oen_psync <= 0;
	else oen_psync <= oen_inv;
always @(negedge clk or posedge rst or negedge set_)
	if(~set_) oen_nsync <= 1;
	else if(rst) oen_nsync <= 0;
	else oen_nsync <= oen_inv;

wire	oen_sel;
assign oen_sel =({CFG_OEN_SEL,init_b} == 5'b00011) ? oen_nsync :
				({CFG_OEN_SEL,init_b} == 5'b00101) ? oen_psync :
				({CFG_OEN_SEL,init_b} == 5'b01001) ? oen_inv:
				({CFG_OEN_SEL,init_b} == 5'b10001) ? 1'b0:
				({CFG_OEN_SEL,init_b} == 5'b00000) ? 1'b1:
				({CFG_OEN_SEL,init_b} == 5'b00001) ? 1'b1 : 1'bx;
assign f_oen = !(gbl_clear_b & ~oen_sel);
endmodule
