module mipi_rx_pinf_tx_pinf_1080 
(
phone_rst,
rx_decode_hsync,
rx_decode_vsync,
swire
);
input phone_rst ;
output rx_decode_hsync ;
output rx_decode_vsync ;
output swire ;
wire phone_rst ;
wire rx_decode_hsync ;
wire rx_decode_vsync ;
wire swire ;
wire \ii2915|xy_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[14]|qx_net  ;
wire \glue_pasm_tx_act_d_reg|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ;
wire \ii2075|xy_net  ;
wire \ii2461|xy_net  ;
wire \ii2846|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21]|qx_net  ;
wire \ii3332|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19]|qx_net  ;
wire \carry_11_ADD_10|s_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[5]|qx_net  ;
wire \ii2777|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2]|qx_net  ;
wire \carry_9_5__ADD_4|co_net  ;
wire \carry_9_8__ADD_7|co_net  ;
wire \ii2333|xy_net  ;
wire \ii2718|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52]|qx_net  ;
wire \carry_12_ADD_10|s_net  ;
wire \carry_12_1__ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[9]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ;
wire \ii2650|xy_net  ;
wire \ii2649|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[10]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[26]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[4]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[21]_net  ;
wire \ii2205|xy_net  ;
wire \ii2195|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8]|qx_net  ;
wire \ii2581|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rstf_reg|qx_net  ;
wire \carry_13_ADD_10|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|almostempty_net  ;
wire \ii2136|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]|qx_net  ;
wire \ii2522|xy_net  ;
wire \ii2897|xy_net  ;
wire \ii2907|xy_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2]|qx_net  ;
wire \ii3383|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ;
wire \ii2067|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg|qx_net  ;
wire \ii2453|xy_net  ;
wire \ii2838|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21]|qx_net  ;
wire \ii3324|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[1]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13]|qx_net  ;
wire \ii2769|xy_net  ;
wire \ii2770|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[21]_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22]|qx_net  ;
wire \carry_9_8__ADD_0|co_net  ;
wire \u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly|xy_net  ;
wire \ii2711|xy_net  ;
wire \carry_9_ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ;
wire \carry_9_11__ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[1]_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[4]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf|xy_net  ;
wire \ii2642|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0]|qx_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3]|qx_net  ;
wire \ii2187|xy_net  ;
wire \ii2573|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13]|qx_net  ;
wire \ii2128|xy_net  ;
wire \ii2514|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7]|qx_net  ;
wire \ii2889|xy_net  ;
wire \ii2890|xy_net  ;
wire \ii2900|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6]|qx_net  ;
wire \ii3375|xy_net  ;
wire \carry_9_3__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_d_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[18]|qx_net  ;
wire \ii2059|xy_net  ;
wire \ii2060|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[27]_net  ;
wire \ii2445|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4]|qx_net  ;
wire \ii2831|xy_net  ;
wire \ii3316|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ;
wire \carry_9_ADD_6|s_net  ;
wire \ii2001|xy_net  ;
wire \ii2376|xy_net  ;
wire \ii2762|xy_net  ;
wire \carry_13_ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0]|qx_net  ;
wire \ii2703|xy_net  ;
wire \ii2693|xy_net  ;
wire \mcu_arbiter_fifo_wr_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6]|qx_net  ;
wire \ii2248|xy_net  ;
wire \ii2634|xy_net  ;
wire \mipi_inst_u_mipi2|CN[0]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[31]|qx_net  ;
wire \ii2179|xy_net  ;
wire \ii2180|xy_net  ;
wire \ii2565|xy_net  ;
wire \ii2121|xy_net  ;
wire \ii2506|xy_net  ;
wire \ii2496|xy_net  ;
wire \ii2882|xy_net  ;
wire \ii3367|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg|qx_net  ;
wire \mcu_arbiter_reg_din_reg[2]|qx_net  ;
wire \carry_9_3__ADD_1|co_net  ;
wire \mipi_inst_u_mipi1|prdata[8]_net  ;
wire \carry_9_6__ADD_4|co_net  ;
wire \carry_9_9__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[5]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1]|qx_net  ;
wire \ii2052|xy_net  ;
wire \ii2437|xy_net  ;
wire \ii2823|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9]|qx_net  ;
wire \ii3308|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2]|qx_net  ;
wire \carry_12_2__ADD_3|co_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[5]_net  ;
wire \carry_13_ADD_8|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3]|qx_net  ;
wire \ii2368|xy_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[1]_net  ;
wire \ii2754|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[17]_net  ;
wire \mipi_inst_u_mipi2|prdata[22]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2]|qx_net  ;
wire \ii2299|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3]|qx_net  ;
wire \ii2685|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[14]_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[22]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[31]_net  ;
wire \carry_8_ADD_3|co_net  ;
wire \ii2241|xy_net  ;
wire \ii2626|xy_net  ;
wire \mcu_arbiter_func_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[14]_net  ;
wire \ii2172|xy_net  ;
wire \ii2557|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0]|qx_net  ;
wire \carry_9_ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9]|qx_net  ;
wire \ii2113|xy_net  ;
wire \ii2488|xy_net  ;
wire \ii2874|xy_net  ;
wire \ii3360|xy_net  ;
wire \ii3359|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[27]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7]|qx_net  ;
wire \carry_11_ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30]|qx_net  ;
wire \carry_9_9__ADD_0|co_net  ;
wire \glue_cmd_s_reg[7]|qx_net  ;
wire \GND_0_inst|Y_net  ;
wire \carry_9_12__ADD_3|co_net  ;
wire \ii2044|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[3]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[3]_net  ;
wire \ii2430|xy_net  ;
wire \ii2429|xy_net  ;
wire \ii2815|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0]|qx_net  ;
wire \ii2746|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11]|qx_net  ;
wire \glue_dnum_s_reg[4]|qx_net  ;
wire \carry_12_ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net  ;
wire \ii2292|xy_net  ;
wire \ii2677|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7]|qx_net  ;
wire \carry_13_ADD_8|co_net  ;
wire \ii2233|xy_net  ;
wire \ii2618|xy_net  ;
wire \carry_9_4__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ;
wire \carry_8_ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0]|qx_net  ;
wire \carry_12_0__ADD_7|co_net  ;
wire \ii2164|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[11]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[9]_net  ;
wire \carry_12_ADD_2|s_net  ;
wire \ii1995|xy_net  ;
wire \ii2095|xy_net  ;
wire \ii2105|xy_net  ;
wire \ii2481|xy_net  ;
wire \ii2866|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23]|qx_net  ;
wire \ii3352|xy_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3]|qx_net  ;
wire \carry_11_ADD_1|co_net  ;
wire \carry_9_10__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22]|qx_net  ;
wire \ii2036|xy_net  ;
wire \ii2422|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[7]|qx_net  ;
wire \ii2797|xy_net  ;
wire \ii2807|xy_net  ;
wire \ii3283|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11]|qx_net  ;
wire \ii2738|xy_net  ;
wire \ii3224|xy_net  ;
wire \carry_12_ADD_1|co_net  ;
wire \mipi_inst_u_mipi2|CM[4]_net  ;
wire \carry_9_11__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[6]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf|xy_net  ;
wire \ii2284|xy_net  ;
wire \ii2670|xy_net  ;
wire \ii2669|xy_net  ;
wire \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|dout[0]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[28]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[5]_net  ;
wire \ii2225|xy_net  ;
wire \carry_13_ADD_1|co_net  ;
wire \ii2611|xy_net  ;
wire \carry_9_4__ADD_1|co_net  ;
wire \carry_9_12__ADD_1|s_net  ;
wire \mipi_inst_u_mipi2|prdata[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2]|qx_net  ;
wire \carry_9_7__ADD_4|co_net  ;
wire \carry_12_ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[10]_net  ;
wire \carry_9_10__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3]|qx_net  ;
wire \carry_12_0__ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[10]_net  ;
wire \ii2156|xy_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[6]_net  ;
wire \ii2927|xy_net  ;
wire \carry_9_10__ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[28]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21]|qx_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[0]_net  ;
wire \carry_9_13__ADD_1|s_net  ;
wire \ii2087|xy_net  ;
wire \ii1987|xy_net  ;
wire \ii2473|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23]|qx_net  ;
wire \ii2858|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[8]_net  ;
wire \ii3344|xy_net  ;
wire \mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[4]_net  ;
wire \carry_9_11__ADD_5|s_net  ;
wire \ii2028|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7]|qx_net  ;
wire \ii2414|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15]|qx_net  ;
wire \ii2789|xy_net  ;
wire \ii2790|xy_net  ;
wire \ii2800|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24]|qx_net  ;
wire \ii2731|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[22]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_valid_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[12]_net  ;
wire \carry_9_12__ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1]|qx_net  ;
wire \ii2662|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5]|qx_net  ;
wire \ii2217|xy_net  ;
wire \ii2603|xy_net  ;
wire \ii2593|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[1]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  ;
wire \carry_9_13__ADD_5|s_net  ;
wire \carry_9_10__ADD_0|co_net  ;
wire \glue_rd_start_s_reg|qx_net  ;
wire \carry_9_13__ADD_3|co_net  ;
wire \mcu_arbiter_u_psram_memack_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15]|qx_net  ;
wire \ii2148|xy_net  ;
wire \ii2919|xy_net  ;
wire \ii2920|xy_net  ;
wire \u_8051_u_h6_8051|memwr_comb_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[21]|qx_net  ;
wire \ii2079|xy_net  ;
wire \ii2080|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6]|qx_net  ;
wire \ii2465|xy_net  ;
wire \ii2851|xy_net  ;
wire \ii3336|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[5]_net  ;
wire \ii2782|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[3]_net  ;
wire \carry_9_5__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1]|qx_net  ;
wire \ii2337|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memack_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2]|qx_net  ;
wire \ii2723|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0]|qx_net  ;
wire \carry_12_1__ADD_7|co_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8]|qx_net  ;
wire \ii2654|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[12]_net  ;
wire \mipi_inst_u_mipi2|prdata[16]_net  ;
wire \ii2199|xy_net  ;
wire \ii2209|xy_net  ;
wire \ii2210|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[11]_net  ;
wire \ii2585|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd_valid_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[8]_net  ;
wire \ii2141|xy_net  ;
wire \ii2526|xy_net  ;
wire \ii2912|xy_net  ;
wire \glue_rx_packet_tx_packet_tx_hsync_fo_reg|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[16]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[25]_net  ;
wire \ii3387|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[29]_net  ;
wire \mipi_inst_u_mipi2|prdata[30]_net  ;
wire \mcu_arbiter_reg_din_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[13]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3]|qx_net  ;
wire \ii2072|xy_net  ;
wire \ii2457|xy_net  ;
wire \ii2843|xy_net  ;
wire \ii3328|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[29]_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[30]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0]|qx_net  ;
wire \carry_11_ADD_4|s_net  ;
wire \ii2774|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[22]_net  ;
wire \carry_9_5__ADD_1|co_net  ;
wire \carry_9_8__ADD_4|co_net  ;
wire \ii2329|xy_net  ;
wire \ii2330|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5]|qx_net  ;
wire \ii2715|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0]|qx_net  ;
wire \carry_9_11__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5]|qx_net  ;
wire \carry_12_1__ADD_0|co_net  ;
wire \ii2646|xy_net  ;
wire \mcu_arbiter_func_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14]|qx_net  ;
wire \carry_12_2__ADD_10|co_net  ;
wire \ii2202|xy_net  ;
wire \ii2192|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[11]_net  ;
wire \ii2577|xy_net  ;
wire \ii2963|xy_net  ;
wire \mcu_arbiter_reg_sel_reg|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi_pll|CLKOUT2_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3]|qx_net  ;
wire \carry_9_3__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1]|qx_net  ;
wire \ii2518|xy_net  ;
wire \ii2894|xy_net  ;
wire \ii2904|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[4]_net  ;
wire \ii3379|xy_net  ;
wire \ii3380|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9]|qx_net  ;
wire \carry_11_ADD_8|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[5]|qx_net  ;
wire \ii2064|xy_net  ;
wire \ii2449|xy_net  ;
wire \ii2450|xy_net  ;
wire \ii2835|xy_net  ;
wire \ii3321|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[6]_net  ;
wire \u_pll_pll_u0|CO2_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2]|qx_net  ;
wire \carry_9_4__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2]|qx_net  ;
wire \ii2381|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13]|qx_net  ;
wire \ii2766|xy_net  ;
wire \glue_dnum_s_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ;
wire \ii2707|xy_net  ;
wire \ii2697|xy_net  ;
wire \carry_9_11__ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3]|qx_net  ;
wire \carry_9_5__ADD_1|s_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net  ;
wire \u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[6]_net  ;
wire \ii2253|xy_net  ;
wire \ii2638|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1]|qx_net  ;
wire \mipi_inst_u_mipi2|host_tx_active_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ;
wire \carry_9_3__ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2]|qx_net  ;
wire \ii2184|xy_net  ;
wire \ii2569|xy_net  ;
wire \ii2570|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf|xy_net  ;
wire \carry_9_6__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[2]_net  ;
wire \glue_rx_packet_tx_packet_tx_vsync_fo_reg|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1]|qx_net  ;
wire \ii2125|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1]|qx_net  ;
wire \ii2511|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[10]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]|qx_net  ;
wire \ii2886|xy_net  ;
wire \carry_9_4__ADD_5|s_net  ;
wire \ii3372|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[0]_net  ;
wire \mipi_inst_u_mipi1|RxActiveHS_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2]|qx_net  ;
wire \carry_9_3__ADD_5|co_net  ;
wire \mipi_inst_u_mipi2|prdata[3]_net  ;
wire \carry_9_6__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24]|qx_net  ;
wire \carry_9_7__ADD_1|s_net  ;
wire \ii2056|xy_net  ;
wire \ii2442|xy_net  ;
wire \ii2827|xy_net  ;
wire \ii3313|xy_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[1]_net  ;
wire \carry_12_2__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[23]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[8]_net  ;
wire \carry_9_5__ADD_5|s_net  ;
wire \ii2373|xy_net  ;
wire \ii2758|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload_valid_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[3]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload_valid_last_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[14]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56]|qx_net  ;
wire \carry_9_8__ADD_1|s_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[6]_net  ;
wire \ii2689|xy_net  ;
wire \ii2690|xy_net  ;
wire \ii2700|xy_net  ;
wire \mcu_arbiter_fifo_clr_f_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf|xy_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[31]|qx_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[7]_net  ;
wire \carry_9_6__ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14]|qx_net  ;
wire \ii2245|xy_net  ;
wire \ii2631|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0]|qx_net  ;
wire \carry_9_9__ADD_1|s_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[16]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5]|qx_net  ;
wire \ii2176|xy_net  ;
wire \ii2562|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|almostempty_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6]|qx_net  ;
wire \carry_9_7__ADD_5|s_net  ;
wire \carry_12_0__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23]|qx_net  ;
wire \carry_9_ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[10]_net  ;
wire \ii2117|xy_net  ;
wire \ii2493|xy_net  ;
wire \ii2503|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[29]_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[30]_net  ;
wire \ii2878|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25]|qx_net  ;
wire \ii3364|xy_net  ;
wire \carry_9_6__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[0]_net  ;
wire \carry_9_9__ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4]|qx_net  ;
wire \carry_9_12__ADD_7|co_net  ;
wire \ii2048|xy_net  ;
wire \mcu_arbiter_fifo_clr_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5]|qx_net  ;
wire \ii2434|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0]|qx_net  ;
wire \ii2819|xy_net  ;
wire \ii2820|xy_net  ;
wire \ii3305|xy_net  ;
wire \carry_9_8__ADD_5|s_net  ;
wire \carry_12_1__ADD_1|s_net  ;
wire \carry_12_2__ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[8]_net  ;
wire \ii2751|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[5]_net  ;
wire \carry_9_9__ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3]|qx_net  ;
wire \ii2296|xy_net  ;
wire \carry_12_2__ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1]|qx_net  ;
wire \ii2682|xy_net  ;
wire \mipi_inst_u_mipi2|CN[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7]|qx_net  ;
wire \carry_8_ADD_0|co_net  ;
wire \ii2237|xy_net  ;
wire \carry_12_0__ADD_5|s_net  ;
wire \ii2623|xy_net  ;
wire \ii3108|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17]|qx_net  ;
wire \ii2168|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1]|qx_net  ;
wire \carry_9_ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2]|qx_net  ;
wire \carry_12_1__ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[23]|qx_net  ;
wire \ii1999|xy_net  ;
wire \ii2099|xy_net  ;
wire \ii2109|xy_net  ;
wire \ii2110|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0]|qx_net  ;
wire \ii2485|xy_net  ;
wire \ii2871|xy_net  ;
wire \ii3356|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3]|qx_net  ;
wire \carry_11_ADD_5|co_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3]|qx_net  ;
wire \carry_9_12__ADD_0|co_net  ;
wire \ii2041|xy_net  ;
wire \ii2426|xy_net  ;
wire \ii2812|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[3]_net  ;
wire \mipi_inst_u_mipi1|pready_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[11]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[19]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[20]_net  ;
wire \carry_12_2__ADD_5|s_net  ;
wire \mipi_inst_u_mipi2|prdata[24]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3]|qx_net  ;
wire \ii2743|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2]|qx_net  ;
wire \carry_12_ADD_5|co_net  ;
wire \glue_rx_packet_tx_packet_rx_active_hs_d_reg|qx_net  ;
wire \carry_12_0__ADD_9|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29]|qx_net  ;
wire \ii2288|xy_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[24]_net  ;
wire \ii2674|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[17]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[16]_net  ;
wire \ii2230|xy_net  ;
wire \ii2229|xy_net  ;
wire \carry_13_ADD_5|co_net  ;
wire \carry_9_4__ADD_5|co_net  ;
wire \ii2615|xy_net  ;
wire \carry_9_7__ADD_8|co_net  ;
wire \carry_12_1__ADD_9|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]|qx_net  ;
wire \carry_12_0__ADD_4|co_net  ;
wire \ii2161|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[11]_net  ;
wire \ii2932|xy_net  ;
wire \mcu_arbiter_reg_din_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[29]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg|qx_net  ;
wire \ii2102|xy_net  ;
wire \ii2092|xy_net  ;
wire \ii1992|xy_net  ;
wire \ii2477|xy_net  ;
wire \carry_12_2__ADD_9|s_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[5]_net  ;
wire \ii2863|xy_net  ;
wire \ii3348|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1]|qx_net  ;
wire \ii2033|xy_net  ;
wire \ii2418|xy_net  ;
wire \ii2804|xy_net  ;
wire \ii2794|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[29]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net  ;
wire \glue_cmd_s_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2]|qx_net  ;
wire \ii2735|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[1]_net  ;
wire \carry_12_0__ADD_10|co_net  ;
wire \ii2281|xy_net  ;
wire \ii2666|xy_net  ;
wire \mcu_arbiter_func_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_tx_cmd_ack_net  ;
wire \ii2222|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[6]_net  ;
wire \ii2607|xy_net  ;
wire \ii2597|xy_net  ;
wire \carry_9_7__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[10]_net  ;
wire \carry_9_10__ADD_4|co_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4]|qx_net  ;
wire \carry_9_13__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0]|qx_net  ;
wire \ii2153|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3]|qx_net  ;
wire \ii2924|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[17]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ;
wire \carry_12_ADD_11|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf|xy_net  ;
wire \ii2084|xy_net  ;
wire \ii1984|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[7]|qx_net  ;
wire \ii2470|xy_net  ;
wire \ii2469|xy_net  ;
wire \ii2855|xy_net  ;
wire \ii3341|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ;
wire \ii2411|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4]|qx_net  ;
wire \ii2786|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15]|qx_net  ;
wire \glue_dnum_s_reg[8]|qx_net  ;
wire \carry_13_ADD_11|s_net  ;
wire \mipi_inst_u_mipi2|CM[6]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[8]_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[9]_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[0]|qx_net  ;
wire \ii2727|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[17]_net  ;
wire \ii2658|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[7]_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg|qx_net  ;
wire \ii2214|xy_net  ;
wire \ii2600|xy_net  ;
wire \ii2590|xy_net  ;
wire \ii2589|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[1]_net  ;
wire \mipi_inst_u_mipi1|prdata[31]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[21]|qx_net  ;
wire \ii1982_dup|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2]|qx_net  ;
wire \carry_9_13__ADD_0|co_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3]|qx_net  ;
wire \ii2145|xy_net  ;
wire \carry_9_ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3]|qx_net  ;
wire \ii2916|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[6]_net  ;
wire \ii2076|xy_net  ;
wire \ii2462|xy_net  ;
wire \ii2847|xy_net  ;
wire \carry_13_ADD_1|s_net  ;
wire \ii3333|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15]|qx_net  ;
wire \ii2778|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[24]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[14]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58]|qx_net  ;
wire \carry_9_5__ADD_5|co_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0]|qx_net  ;
wire \carry_9_8__ADD_8|co_net  ;
wire \ii2334|xy_net  ;
wire \ii2720|xy_net  ;
wire \ii2719|xy_net  ;
wire \ii3195|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3]|qx_net  ;
wire \carry_12_1__ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16]|qx_net  ;
wire \ii2651|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[3]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[7]_net  ;
wire \carry_9_ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7]|qx_net  ;
wire \ii2206|xy_net  ;
wire \ii2196|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[5]_net  ;
wire \ii2582|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_valid_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25]|qx_net  ;
wire \carry_13_ADD_5|s_net  ;
wire \ii2137|xy_net  ;
wire \ii2523|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27]|qx_net  ;
wire \ii2908|xy_net  ;
wire \ii2898|xy_net  ;
wire \ii3384|xy_net  ;
wire \carry_12_0__ADD_10|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7]|qx_net  ;
wire \ii2068|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[7]_net  ;
wire \ii2454|xy_net  ;
wire \ii2840|xy_net  ;
wire \ii2839|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0]|qx_net  ;
wire \ii3325|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_d_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[5]_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28]|qx_net  ;
wire \ii2771|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[2]_net  ;
wire \carry_9_8__ADD_1|co_net  ;
wire \ii2712|xy_net  ;
wire \carry_9_11__ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[14]_net  ;
wire \mipi_inst_u_mipi2|prdata[18]_net  ;
wire \ii2643|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ;
wire \carry_13_ADD_9|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1]|qx_net  ;
wire \ii2188|xy_net  ;
wire \ii2574|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[27]_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[18]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[25]|qx_net  ;
wire \ii2129|xy_net  ;
wire \ii2130|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]|qx_net  ;
wire \ii2515|xy_net  ;
wire \ii2891|xy_net  ;
wire \ii2901|xy_net  ;
wire \ii3376|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5]|qx_net  ;
wire \ii2061|xy_net  ;
wire \ii2446|xy_net  ;
wire \ii2832|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4]|qx_net  ;
wire \ii3317|xy_net  ;
wire \mipi_inst_u_mipi2|host_tx_payload_en_last_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[24]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7]|qx_net  ;
wire \ii2377|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6]|qx_net  ;
wire \ii2763|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[0]_net  ;
wire \mipi_inst_u_mipi_pll|LOCK_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16]|qx_net  ;
wire \carry_8_ADD_1|s_net  ;
wire \ii2704|xy_net  ;
wire \ii2694|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[19]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12]|qx_net  ;
wire \glue_dnum_s_reg[11]|qx_net  ;
wire \u_8051_u_h6_8051|mempsrd_comb_net  ;
wire \u_8051_u_h6_8051|port0o[0]_net  ;
wire \ii2249|xy_net  ;
wire \ii2250|xy_net  ;
wire \u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly|xy_net  ;
wire \ii2635|xy_net  ;
wire \mipi_inst_u_mipi2|CO[0]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]|qx_net  ;
wire \ii2181|xy_net  ;
wire \ii2566|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[8]|qx_net  ;
wire \ii2122|xy_net  ;
wire \ii2507|xy_net  ;
wire \ii2497|xy_net  ;
wire \VCC_0_inst|Y_net  ;
wire \ii2883|xy_net  ;
wire \ii3368|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net  ;
wire \carry_9_3__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[8]_net  ;
wire \carry_9_6__ADD_5|co_net  ;
wire \carry_9_9__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3]|qx_net  ;
wire \ii2053|xy_net  ;
wire \ii2438|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[6]_net  ;
wire \ii2824|xy_net  ;
wire \ii3310|xy_net  ;
wire \ii3309|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3]|qx_net  ;
wire \carry_12_2__ADD_4|co_net  ;
wire \carry_8_ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_dphy_direction_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[12]_net  ;
wire \glue_cmd_s_reg[2]|qx_net  ;
wire \ii2369|xy_net  ;
wire \ii2370|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net  ;
wire \ii2755|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[14]_net  ;
wire \carry_12_ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[8]_net  ;
wire \ii2686|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1]|qx_net  ;
wire \carry_9_10__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18]|qx_net  ;
wire \mipi_inst_u_mipi2|CM[1]_net  ;
wire \carry_12_1__ADD_10|s_net  ;
wire \ii2242|xy_net  ;
wire \carry_8_ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0]|qx_net  ;
wire \ii2627|xy_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2]|qx_net  ;
wire \ii2173|xy_net  ;
wire \ii2558|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[12]_net  ;
wire \carry_9_11__ADD_2|s_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[5]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[10]_net  ;
wire \carry_9_ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[9]|qx_net  ;
wire \ii2114|xy_net  ;
wire \ii2489|xy_net  ;
wire \ii2490|xy_net  ;
wire \ii2500|xy_net  ;
wire \ii2875|xy_net  ;
wire \ii3361|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[11]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[3]_net  ;
wire \carry_11_ADD_9|co_net  ;
wire \carry_9_9__ADD_1|co_net  ;
wire \mipi_inst_u_mipi1|prdata[25]_net  ;
wire \carry_9_12__ADD_4|co_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf|xy_net  ;
wire \ii2045|xy_net  ;
wire \carry_9_12__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6]|qx_net  ;
wire \ii2431|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17]|qx_net  ;
wire \carry_12_ADD_7|s_net  ;
wire \ii2816|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[8]_net  ;
wire \carry_9_10__ADD_6|s_net  ;
wire \ii2747|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[1]_net  ;
wire \carry_12_ADD_9|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2]|qx_net  ;
wire \carry_9_13__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4]|qx_net  ;
wire \ii2293|xy_net  ;
wire \ii2678|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[18]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6]|qx_net  ;
wire \carry_9_11__ADD_6|s_net  ;
wire \ii2234|xy_net  ;
wire \carry_13_ADD_9|co_net  ;
wire \ii2619|xy_net  ;
wire \ii2620|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[23]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0]|qx_net  ;
wire \carry_12_0__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  ;
wire \ii2165|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6]|qx_net  ;
wire \carry_9_12__ADD_6|s_net  ;
wire \u_pll_pll_u0|CO0_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]|qx_net  ;
wire \ii2106|xy_net  ;
wire \ii2096|xy_net  ;
wire \ii1996|xy_net  ;
wire \ii2482|xy_net  ;
wire \ii2867|xy_net  ;
wire \ii3353|xy_net  ;
wire \carry_11_ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15]|qx_net  ;
wire \ii2037|xy_net  ;
wire \ii2423|xy_net  ;
wire \ii2808|xy_net  ;
wire \ii2798|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17]|qx_net  ;
wire \ii3284|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[7]_net  ;
wire \carry_9_13__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10]|qx_net  ;
wire \ii2739|xy_net  ;
wire \ii2740|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5]|qx_net  ;
wire \carry_12_ADD_2|co_net  ;
wire \mipi_inst_u_mipi2|CN[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18]|qx_net  ;
wire \ii2285|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[0]_net  ;
wire \ii2671|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1]|qx_net  ;
wire \carry_13_ADD_2|co_net  ;
wire \ii2226|xy_net  ;
wire \carry_9_4__ADD_2|co_net  ;
wire \ii2612|xy_net  ;
wire \carry_9_7__ADD_5|co_net  ;
wire \carry_9_10__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[11]_net  ;
wire \carry_12_0__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[9]_net  ;
wire \ii2157|xy_net  ;
wire \ii2928|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[13]_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30]|qx_net  ;
wire \carry_11_ADD_1|s_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2]|qx_net  ;
wire \ii1988|xy_net  ;
wire \ii2088|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9]|qx_net  ;
wire \ii2474|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4]|qx_net  ;
wire \ii2859|xy_net  ;
wire \ii2860|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3]|qx_net  ;
wire \ii3345|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[5]_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_d_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[22]_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[13]_net  ;
wire \mipi_inst_u_mipi2|prdata[26]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[10]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31]|qx_net  ;
wire \ii2030|xy_net  ;
wire \ii2029|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1]|qx_net  ;
wire \ii2415|xy_net  ;
wire \ii2801|xy_net  ;
wire \ii2791|xy_net  ;
wire \carry_12_2__ADD_10|s_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[26]_net  ;
wire \ii2732|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6]|qx_net  ;
wire \u_pll_pll_u0|PLOCK_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[18]_net  ;
wire \ii2663|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3]|qx_net  ;
wire \carry_11_ADD_5|s_net  ;
wire \ii2218|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ;
wire \ii2594|xy_net  ;
wire \ii2604|xy_net  ;
wire \ii3079|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net  ;
wire \carry_9_10__ADD_1|co_net  ;
wire \carry_9_13__ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6]|qx_net  ;
wire \ii2150|xy_net  ;
wire \ii2149|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[27]|qx_net  ;
wire \ii3021|xy_net  ;
wire \ii2921|xy_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7]|qx_net  ;
wire \ii2081|xy_net  ;
wire \ii2466|xy_net  ;
wire \ii2852|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net  ;
wire \ii3337|xy_net  ;
wire \rstn_r_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_fifo_readen_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7]|qx_net  ;
wire \ii2783|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[3]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18]|qx_net  ;
wire \carry_9_3__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0]|qx_net  ;
wire \ii2338|xy_net  ;
wire \ii2724|xy_net  ;
wire \mcu_arbiter_data_sel_reg|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[22]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6]|qx_net  ;
wire \carry_11_ADD_9|s_net  ;
wire \glue_dnum_s_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14]|qx_net  ;
wire \carry_12_1__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0]|qx_net  ;
wire \ii2655|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0]|qx_net  ;
wire \carry_9_4__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_rstsf_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  ;
wire \ii2211|xy_net  ;
wire \ii2586|xy_net  ;
wire \mcu_arbiter_func_reg[0]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[19]_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[20]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3]|qx_net  ;
wire \ii2142|xy_net  ;
wire \ii2913|xy_net  ;
wire \ii3388|xy_net  ;
wire \carry_9_5__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5]|qx_net  ;
wire \ii2073|xy_net  ;
wire \ii2458|xy_net  ;
wire \ii2844|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf|xy_net  ;
wire \ii3329|xy_net  ;
wire \ii3330|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3]|qx_net  ;
wire \carry_9_3__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[0]_net  ;
wire \glue_cmd_s_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[0]|qx_net  ;
wire \carry_9_6__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6]|qx_net  ;
wire \ii2775|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ;
wire \carry_9_5__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  ;
wire \carry_9_8__ADD_5|co_net  ;
wire \mipi_inst_u_mipi1|prdata[20]_net  ;
wire \mipi_inst_u_mipi1|prdata[19]_net  ;
wire \ii2331|xy_net  ;
wire \ii2716|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[5]_net  ;
wire \carry_9_4__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[9]_net  ;
wire \carry_9_11__ADD_8|co_net  ;
wire \glue_dnum_s_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5]|qx_net  ;
wire \carry_12_1__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21]|qx_net  ;
wire \carry_9_7__ADD_2|s_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[11]_net  ;
wire \ii2647|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[3]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3]|qx_net  ;
wire \io_phone_rst_inst|f_id[0]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23]|qx_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[4]_net  ;
wire \carry_9_5__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4]|qx_net  ;
wire \ii2193|xy_net  ;
wire \ii2203|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7]|qx_net  ;
wire \ii2578|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ;
wire \carry_9_8__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[13]_net  ;
wire \ii2134|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[8]_net  ;
wire \ii2520|xy_net  ;
wire \ii2519|xy_net  ;
wire \ii2905|xy_net  ;
wire \ii2895|xy_net  ;
wire \ii3381|xy_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[13]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ;
wire \carry_9_6__ADD_6|s_net  ;
wire \ii2065|xy_net  ;
wire \ii2451|xy_net  ;
wire \ii2836|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20]|qx_net  ;
wire \ii3322|xy_net  ;
wire \carry_9_9__ADD_2|s_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[26]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18]|qx_net  ;
wire \ii2767|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[4]|qx_net  ;
wire \ii3253|xy_net  ;
wire \carry_9_7__ADD_6|s_net  ;
wire \carry_12_0__ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1]|qx_net  ;
wire \ii2698|xy_net  ;
wire \ii2708|xy_net  ;
wire \carry_9_11__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[5]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1]|qx_net  ;
wire \ii2254|xy_net  ;
wire \ii2640|xy_net  ;
wire \ii2639|xy_net  ;
wire \carry_9_8__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5]|qx_net  ;
wire \carry_12_1__ADD_2|s_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_frame_start_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7]|qx_net  ;
wire \ii2185|xy_net  ;
wire \ii2571|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0]|qx_net  ;
wire \carry_9_9__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31]|qx_net  ;
wire \carry_12_2__ADD_2|s_net  ;
wire \ii2126|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]|qx_net  ;
wire \ii2512|xy_net  ;
wire \ii2887|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1]|qx_net  ;
wire \ii3373|xy_net  ;
wire \carry_9_3__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[7]_net  ;
wire \ii2057|xy_net  ;
wire \carry_12_0__ADD_6|s_net  ;
wire \ii2443|xy_net  ;
wire \ii2828|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20]|qx_net  ;
wire \ii3314|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[4]_net  ;
wire \carry_12_2__ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12]|qx_net  ;
wire \ii2374|xy_net  ;
wire \ii2760|xy_net  ;
wire \ii2759|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13]|qx_net  ;
wire \carry_12_1__ADD_6|s_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[16]_net  ;
wire \mipi_inst_u_mipi2|prdata[21]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21]|qx_net  ;
wire \ii2701|xy_net  ;
wire \ii2691|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3]|qx_net  ;
wire \ii2246|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[13]_net  ;
wire \ii2632|xy_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[21]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[29]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[30]_net  ;
wire \carry_12_2__ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]|qx_net  ;
wire \ii2177|xy_net  ;
wire \ii2563|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[6]_net  ;
wire \mcu_arbiter_u_emif2apb_memrd_s_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12]|qx_net  ;
wire \carry_9_ADD_8|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4]|qx_net  ;
wire \ii2118|xy_net  ;
wire \ii2504|xy_net  ;
wire \ii2494|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4]|qx_net  ;
wire \ii2880|xy_net  ;
wire \ii2879|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4]|qx_net  ;
wire \ii3365|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5]|qx_net  ;
wire \carry_9_6__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_d_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5]|qx_net  ;
wire \carry_9_9__ADD_5|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[26]_net  ;
wire \carry_9_12__ADD_8|co_net  ;
wire \ii2050|xy_net  ;
wire \ii2049|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[17]|qx_net  ;
wire \ii2435|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3]|qx_net  ;
wire \ii2821|xy_net  ;
wire \ii3306|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ;
wire \carry_12_2__ADD_1|co_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[2]_net  ;
wire \ii2752|xy_net  ;
wire \ii2297|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0]|qx_net  ;
wire \ii2683|xy_net  ;
wire \u_8051_u_h6_8051|port0o[2]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5]|qx_net  ;
wire \ii2238|xy_net  ;
wire \carry_8_ADD_1|co_net  ;
wire \ii2624|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[12]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[8]_net  ;
wire \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net  ;
wire \ii2170|xy_net  ;
wire \ii2169|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[30]|qx_net  ;
wire \ii2555|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[10]_net  ;
wire \carry_9_ADD_1|co_net  ;
wire \ii2111|xy_net  ;
wire \ii2486|xy_net  ;
wire \ii2872|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[8]_net  ;
wire \ii3357|xy_net  ;
wire \mcu_arbiter_reg_din_reg[1]|qx_net  ;
wire \carry_11_ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[14]_net  ;
wire \carry_9_12__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[1]|qx_net  ;
wire \ii2042|xy_net  ;
wire \ii2427|xy_net  ;
wire \ii2813|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[15]_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2]|qx_net  ;
wire \ii2744|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf|xy_net  ;
wire \carry_12_ADD_6|co_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8]|qx_net  ;
wire \glue_dnum_s_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0]|qx_net  ;
wire \mipi_inst_u_mipi2|host_tx_payload_en_net  ;
wire \mipi_inst_u_mipi2|CM[3]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1]|qx_net  ;
wire \ii2300|xy_net  ;
wire \ii2290|xy_net  ;
wire \ii2289|xy_net  ;
wire \ii2675|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[5]_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[6]_net  ;
wire \carry_9_ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf|xy_net  ;
wire \ii2231|xy_net  ;
wire \carry_13_ADD_6|co_net  ;
wire \carry_9_4__ADD_6|co_net  ;
wire \ii2616|xy_net  ;
wire \ii2992|xy_net  ;
wire \carry_13_ADD_12|s_net  ;
wire \mcu_arbiter_func_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[4]_net  ;
wire \mipi_inst_u_mipi2|prdata[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  ;
wire \carry_12_0__ADD_5|co_net  ;
wire \ii2162|xy_net  ;
wire \ii2933|xy_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[5]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[27]_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11]|qx_net  ;
wire \ii2103|xy_net  ;
wire \ii2093|xy_net  ;
wire \ii1993|xy_net  ;
wire \ii2478|xy_net  ;
wire \ii2864|xy_net  ;
wire \ii3350|xy_net  ;
wire \ii3349|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[7]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28]|qx_net  ;
wire \glue_cmd_s_reg[6]|qx_net  ;
wire \ii2034|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[2]|qx_net  ;
wire \ii2420|xy_net  ;
wire \ii2419|xy_net  ;
wire \ii2805|xy_net  ;
wire \ii2795|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[3]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12]|qx_net  ;
wire \carry_9_ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ;
wire \ii2736|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10]|qx_net  ;
wire \glue_dnum_s_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[21]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[11]_net  ;
wire \ii2282|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4]|qx_net  ;
wire \carry_13_ADD_2|s_net  ;
wire \ii2667|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6]|qx_net  ;
wire \ii2223|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ;
wire \ii2608|xy_net  ;
wire \ii2598|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1]|qx_net  ;
wire \carry_9_7__ADD_2|co_net  ;
wire \carry_9_10__ADD_5|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41]|qx_net  ;
wire \carry_9_13__ADD_8|co_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[11]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[4]_net  ;
wire \ii2154|xy_net  ;
wire \ii2925|xy_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg|qx_net  ;
wire \ii2085|xy_net  ;
wire \ii1985|xy_net  ;
wire \ii2471|xy_net  ;
wire \ii2856|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22]|qx_net  ;
wire \ii3342|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0]|qx_net  ;
wire \u_osc|OSC_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21]|qx_net  ;
wire \ii2026|xy_net  ;
wire \ii2412|xy_net  ;
wire \ii2787|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6]|qx_net  ;
wire \carry_13_ADD_6|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10]|qx_net  ;
wire \ii2728|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[2]_net  ;
wire \carry_12_0__ADD_11|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t105_out1_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3]|qx_net  ;
wire \ii2660|xy_net  ;
wire \ii2659|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ;
wire \ii2215|xy_net  ;
wire \ii2601|xy_net  ;
wire \ii2591|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[10]_net  ;
wire \carry_9_13__ADD_1|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]|qx_net  ;
wire \ii2146|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]|qx_net  ;
wire \ii2917|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[15]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[24]_net  ;
wire \mipi_inst_u_mipi2|prdata[28]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[12]_net  ;
wire \ii2077|xy_net  ;
wire \ii2463|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22]|qx_net  ;
wire \ii2848|xy_net  ;
wire \ii3334|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14]|qx_net  ;
wire \ii2780|xy_net  ;
wire \ii2779|xy_net  ;
wire \u_pll_pll_u0|CO3_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[28]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15]|qx_net  ;
wire \carry_9_5__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23]|qx_net  ;
wire \ii2335|xy_net  ;
wire \glue_rx_packet_tx_packet_fifo_vs_reg|qx_net  ;
wire \ii2721|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[21]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8]|qx_net  ;
wire \carry_12_1__ADD_5|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0]|qx_net  ;
wire \ii2652|xy_net  ;
wire \ii3137|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  ;
wire \ii2207|xy_net  ;
wire \ii2197|xy_net  ;
wire \ii2583|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[9]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14]|qx_net  ;
wire \carry_8_ADD_2|s_net  ;
wire \ii2138|xy_net  ;
wire \ii2524|xy_net  ;
wire \ii2910|xy_net  ;
wire \ii2909|xy_net  ;
wire \ii2899|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6]|qx_net  ;
wire \ii3385|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7]|qx_net  ;
wire \ii2070|xy_net  ;
wire \ii2069|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[20]|qx_net  ;
wire \mcu_arbiter_mipi_sel_reg|qx_net  ;
wire \ii2455|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5]|qx_net  ;
wire \ii2841|xy_net  ;
wire \ii3326|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0]|qx_net  ;
wire \ii2772|xy_net  ;
wire \glue_rx_packet_tx_packet_sc_vs_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0]|qx_net  ;
wire \u_8051_u_h6_8051|mempswr_comb_net  ;
wire \carry_9_8__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0]|qx_net  ;
wire \ii2713|xy_net  ;
wire \carry_9_11__ADD_5|co_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ;
wire \ii2644|xy_net  ;
wire \carry_8_ADD_6|s_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[5]_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[22]_net  ;
wire \ii2200|xy_net  ;
wire \ii2190|xy_net  ;
wire \ii2189|xy_net  ;
wire \ii2575|xy_net  ;
wire \carry_12_ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[1]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t71_out1_reg|qx_net  ;
wire \ii2131|xy_net  ;
wire \ii2516|xy_net  ;
wire \ii2892|xy_net  ;
wire \ii2902|xy_net  ;
wire \ii3377|xy_net  ;
wire \carry_9_10__ADD_3|s_net  ;
wire \mcu_arbiter_reg_din_reg[3]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[3]|qx_net  ;
wire \carry_12_1__ADD_11|s_net  ;
wire \ii2062|xy_net  ;
wire \ii2447|xy_net  ;
wire \ii2833|xy_net  ;
wire \ii3318|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4]|qx_net  ;
wire \ii2378|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[22]_net  ;
wire \carry_9_11__ADD_3|s_net  ;
wire \ii2764|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[7]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[26]|qx_net  ;
wire \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[13]_net  ;
wire \ii2705|xy_net  ;
wire \ii2695|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4]|qx_net  ;
wire \mcu_arbiter_apb_sel_reg|qx_net  ;
wire \carry_9_12__ADD_3|s_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[6]_net  ;
wire \ii2251|xy_net  ;
wire \carry_12_ADD_8|s_net  ;
wire \ii2636|xy_net  ;
wire \mcu_arbiter_func_reg[4]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13]|qx_net  ;
wire \carry_9_10__ADD_7|s_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[15]_net  ;
wire \mcu_arbiter_fifo_clr_s_reg|qx_net  ;
wire \ii2182|xy_net  ;
wire \ii2567|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1]|qx_net  ;
wire \carry_9_13__ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi1|tx_dphy_rdy_net  ;
wire \ii2123|xy_net  ;
wire \ii2508|xy_net  ;
wire \ii2498|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0]|qx_net  ;
wire \ii2884|xy_net  ;
wire \ii3370|xy_net  ;
wire \ii3369|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7]|qx_net  ;
wire \carry_9_3__ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8]|qx_net  ;
wire \carry_9_6__ADD_6|co_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[28]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31]|qx_net  ;
wire \carry_9_11__ADD_7|s_net  ;
wire \ii2054|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[4]|qx_net  ;
wire \ii2440|xy_net  ;
wire \ii2439|xy_net  ;
wire \ii2825|xy_net  ;
wire \ii3311|xy_net  ;
wire \carry_12_2__ADD_5|co_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14]|qx_net  ;
wire \ii2371|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1]|qx_net  ;
wire \ii2756|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12]|qx_net  ;
wire \glue_dnum_s_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7]|qx_net  ;
wire \carry_9_12__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11]|qx_net  ;
wire \carry_12_ADD_10|co_net  ;
wire \ii2687|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7]|qx_net  ;
wire \mipi_inst_u_mipi2|CN[1]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27]|qx_net  ;
wire \ii2243|xy_net  ;
wire \carry_8_ADD_5|co_net  ;
wire \ii2628|xy_net  ;
wire \carry_9_13__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ;
wire \ii2174|xy_net  ;
wire \ii2560|xy_net  ;
wire \ii2559|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[17]|qx_net  ;
wire \carry_9_ADD_5|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0]|qx_net  ;
wire \ii2115|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[9]_net  ;
wire \ii2491|xy_net  ;
wire \ii2501|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ;
wire \ii2876|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]|qx_net  ;
wire \ii3362|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[10]_net  ;
wire \carry_9_9__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2]|qx_net  ;
wire \carry_9_12__ADD_5|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[6]_net  ;
wire \ii2046|xy_net  ;
wire \ii2432|xy_net  ;
wire \ii2817|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[10]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[18]_net  ;
wire \mipi_inst_u_mipi2|prdata[23]_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12]|qx_net  ;
wire \ii2748|xy_net  ;
wire \carry_11_ADD_2|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5]|qx_net  ;
wire \ii2294|xy_net  ;
wire \ii2680|xy_net  ;
wire \ii2679|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[15]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[30]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[29]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[23]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13]|qx_net  ;
wire \ii2235|xy_net  ;
wire \ii2621|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[15]_net  ;
wire \carry_12_2__ADD_11|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4]|qx_net  ;
wire \carry_12_0__ADD_9|co_net  ;
wire \ii2166|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[28]_net  ;
wire \ii2107|xy_net  ;
wire \ii2097|xy_net  ;
wire \ii1997|xy_net  ;
wire \ii2483|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24]|qx_net  ;
wire \ii2868|xy_net  ;
wire \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|empty_net  ;
wire \ii3354|xy_net  ;
wire \carry_11_ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[4]_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11]|qx_net  ;
wire \carry_11_ADD_6|s_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4]|qx_net  ;
wire \ii2038|xy_net  ;
wire \ii2424|xy_net  ;
wire \ii2810|xy_net  ;
wire \ii2809|xy_net  ;
wire \ii2799|xy_net  ;
wire \ii3285|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25]|qx_net  ;
wire \ii2741|xy_net  ;
wire \carry_12_ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2]|qx_net  ;
wire \ii2286|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0]|qx_net  ;
wire \ii2672|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6]|qx_net  ;
wire \carry_13_ADD_3|co_net  ;
wire \ii2227|xy_net  ;
wire \carry_9_4__ADD_3|co_net  ;
wire \ii2613|xy_net  ;
wire \carry_9_7__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  ;
wire \carry_9_3__ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16]|qx_net  ;
wire \carry_12_0__ADD_2|co_net  ;
wire \ii2158|xy_net  ;
wire \ii2930|xy_net  ;
wire \ii2929|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0]|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[16]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[22]|qx_net  ;
wire \ii1989|xy_net  ;
wire \ii1990|xy_net  ;
wire \ii2089|xy_net  ;
wire \ii2090|xy_net  ;
wire \ii2100|xy_net  ;
wire \ii2475|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7]|qx_net  ;
wire \ii2861|xy_net  ;
wire \ii3346|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2]|qx_net  ;
wire \carry_9_4__ADD_3|s_net  ;
wire \carry_13_ADD_10|co_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2]|qx_net  ;
wire \ii2031|xy_net  ;
wire \ii2416|xy_net  ;
wire \ii2802|xy_net  ;
wire \ii2792|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi2|CM[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3]|qx_net  ;
wire \ii2733|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1]|qx_net  ;
wire \carry_9_5__ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[7]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|dout[1]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9]|qx_net  ;
wire \ii2664|xy_net  ;
wire \carry_9_3__ADD_7|s_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[16]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[16]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[6]_net  ;
wire \mipi_inst_u_mipi2|prdata[9]_net  ;
wire \carry_9_6__ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[11]_net  ;
wire \ii2219|xy_net  ;
wire \ii2220|xy_net  ;
wire \ii2595|xy_net  ;
wire \ii2605|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ;
wire \carry_9_10__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[11]_net  ;
wire \carry_9_13__ADD_5|co_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[0]_net  ;
wire \mipi_inst_u_mipi1|prdata[29]_net  ;
wire \mipi_inst_u_mipi1|prdata[30]_net  ;
wire \carry_9_4__ADD_7|s_net  ;
wire \ii2151|xy_net  ;
wire \ii2922|xy_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[1]_net  ;
wire \mcu_arbiter_reg_din_reg[5]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[9]_net  ;
wire \carry_9_7__ADD_3|s_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4]|qx_net  ;
wire \ii2082|xy_net  ;
wire \ii1982|xy_net  ;
wire \ii2467|xy_net  ;
wire \ii2853|xy_net  ;
wire \ii3338|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[5]_net  ;
wire \glue_rx_packet_tx_packet_fifo_empty_reg|qx_net  ;
wire \carry_9_5__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0]|qx_net  ;
wire \ii2784|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[28]|qx_net  ;
wire \carry_9_8__ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[23]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[13]_net  ;
wire \ii2339|xy_net  ;
wire \ii2340|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5]|qx_net  ;
wire \ii2725|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2]|qx_net  ;
wire \carry_9_6__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6]|qx_net  ;
wire \carry_12_1__ADD_9|co_net  ;
wire \glue_rd_start_f_reg|qx_net  ;
wire \ii2656|xy_net  ;
wire \carry_9_9__ADD_3|s_net  ;
wire \mcu_arbiter_func_reg[6]|qx_net  ;
wire \carry_12_1__ADD_10|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[2]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[6]_net  ;
wire \ii2212|xy_net  ;
wire \ii2587|xy_net  ;
wire \carry_9_7__ADD_7|s_net  ;
wire \carry_12_0__ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[4]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17]|qx_net  ;
wire \mipi_inst_u_mipi2|tx_dphy_rdy_net  ;
wire \ii2143|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2]|qx_net  ;
wire \ii2914|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ;
wire \glue_pasm_cmd_rq_o_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[6]|qx_net  ;
wire \ii2074|xy_net  ;
wire \carry_9_8__ADD_7|s_net  ;
wire \carry_12_1__ADD_3|s_net  ;
wire \ii2459|xy_net  ;
wire \ii2460|xy_net  ;
wire \ii2845|xy_net  ;
wire \ii3331|xy_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_rd_start_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14]|qx_net  ;
wire \ii2776|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[4]_net  ;
wire \glue_dnum_s_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27]|qx_net  ;
wire \carry_9_9__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2]|qx_net  ;
wire \carry_12_2__ADD_3|s_net  ;
wire \carry_9_5__ADD_3|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1]|qx_net  ;
wire \carry_9_8__ADD_6|co_net  ;
wire \mipi_inst_u_mipi2|pready_net  ;
wire \ii2332|xy_net  ;
wire \ii2717|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[1]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4]|qx_net  ;
wire \carry_12_1__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29]|qx_net  ;
wire \carry_12_0__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ;
wire \ii2648|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[17]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3]|qx_net  ;
wire \ii2194|xy_net  ;
wire \ii2204|xy_net  ;
wire \ii2579|xy_net  ;
wire \ii2580|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[8]_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[20]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[9]_net  ;
wire \carry_12_1__ADD_7|s_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[26]_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[17]_net  ;
wire \mipi_inst_u_mipi2|prdata[31]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[14]_net  ;
wire \ii2135|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2]|qx_net  ;
wire \ii2521|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]|qx_net  ;
wire \ii2906|xy_net  ;
wire \ii2896|xy_net  ;
wire \ii3382|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25]|qx_net  ;
wire \ii2066|xy_net  ;
wire \ii2452|xy_net  ;
wire \ii2837|xy_net  ;
wire \ii3323|xy_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[31]_net  ;
wire \carry_12_2__ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12]|qx_net  ;
wire \ii2768|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[23]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7]|qx_net  ;
wire \ii2710|xy_net  ;
wire \ii2709|xy_net  ;
wire \ii2699|xy_net  ;
wire \carry_9_11__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15]|qx_net  ;
wire \ii2641|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6]|qx_net  ;
wire \ii2186|xy_net  ;
wire \ii2572|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7]|qx_net  ;
wire \u_gbuf_u_gbuf|out_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[5]_net  ;
wire \ii2127|xy_net  ;
wire \ii2513|xy_net  ;
wire \mcu_arbiter_u_emif2apb_fpga_HRD_reg|qx_net  ;
wire \ii2888|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26]|qx_net  ;
wire \ii3374|xy_net  ;
wire \carry_9_3__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[7]_net  ;
wire \ii2058|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6]|qx_net  ;
wire \ii2444|xy_net  ;
wire \ii2830|xy_net  ;
wire \ii2829|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0]|qx_net  ;
wire \ii3315|xy_net  ;
wire \carry_12_2__ADD_9|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[5]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[12]|qx_net  ;
wire \ii2000|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27]|qx_net  ;
wire \ii2375|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[11]_net  ;
wire \ii2761|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[12]_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[13]_net  ;
wire \ii2692|xy_net  ;
wire \ii2702|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8]|qx_net  ;
wire \ii2247|xy_net  ;
wire \ii2633|xy_net  ;
wire \mipi_inst_u_mipi2|CM[0]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2]|qx_net  ;
wire \mipi_inst_u_mipi_pll|CLKOUT1_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[3]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0]|qx_net  ;
wire \ii2178|xy_net  ;
wire \ii2564|xy_net  ;
wire \ii3050|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[1]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[24]|qx_net  ;
wire \ii2119|xy_net  ;
wire \ii2120|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1]|qx_net  ;
wire \ii2495|xy_net  ;
wire \ii2505|xy_net  ;
wire \ii2881|xy_net  ;
wire \ii3366|xy_net  ;
wire \carry_9_ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4]|qx_net  ;
wire \carry_9_3__ADD_0|co_net  ;
wire \u_pll_pll_u0|CO1_net  ;
wire \carry_9_6__ADD_3|co_net  ;
wire \carry_9_9__ADD_6|co_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[2]_net  ;
wire \ii2051|xy_net  ;
wire \ii2436|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2]|qx_net  ;
wire \ii2822|xy_net  ;
wire \mipi_inst_u_mipi1|prdata[24]_net  ;
wire \ii3307|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[9]_net  ;
wire \carry_12_2__ADD_2|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5]|qx_net  ;
wire \ii2753|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[15]_net  ;
wire \mipi_inst_u_mipi2|clk_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[0]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31]|qx_net  ;
wire \ii2298|xy_net  ;
wire \ii2684|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[18]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11]|qx_net  ;
wire \glue_dnum_s_reg[10]|qx_net  ;
wire \carry_8_ADD_2|co_net  ;
wire \ii2239|xy_net  ;
wire \ii2240|xy_net  ;
wire \ii2625|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[17]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]|qx_net  ;
wire \carry_9_ADD_5|s_net  ;
wire \ii2171|xy_net  ;
wire \ii2556|xy_net  ;
wire \mcu_arbiter_reg_din_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[31]_net  ;
wire \carry_9_ADD_2|co_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[7]|qx_net  ;
wire \carry_13_ADD_3|s_net  ;
wire \ii2112|xy_net  ;
wire \ii2487|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[1]_net  ;
wire \ii2873|xy_net  ;
wire \ii3358|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7]|qx_net  ;
wire \carry_11_ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2]|qx_net  ;
wire \carry_9_12__ADD_2|co_net  ;
wire \ii2043|xy_net  ;
wire \ii2428|xy_net  ;
wire \ii2814|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_cmd_s_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7]|qx_net  ;
wire \ii2745|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8]|qx_net  ;
wire \carry_12_ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0]|qx_net  ;
wire \mipi_inst_u_mipi2|CN[3]_net  ;
wire \ii2291|xy_net  ;
wire \ii2301|xy_net  ;
wire \ii2676|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0]|qx_net  ;
wire \glue_pasm_packet_finish_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17]|qx_net  ;
wire \carry_13_ADD_7|co_net  ;
wire \ii2232|xy_net  ;
wire \ii2617|xy_net  ;
wire \carry_9_4__ADD_7|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5]|qx_net  ;
wire \carry_13_ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6]|qx_net  ;
wire \carry_12_0__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1]|qx_net  ;
wire \ii2163|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4]|qx_net  ;
wire \ii2934|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[8]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[12]_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[8]|qx_net  ;
wire \ii1994|xy_net  ;
wire \ii2094|xy_net  ;
wire \ii2104|xy_net  ;
wire \ii2479|xy_net  ;
wire \ii2480|xy_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[8]_net  ;
wire \ii2865|xy_net  ;
wire \ii3351|xy_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[10]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5]|qx_net  ;
wire \carry_11_ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[4]_net  ;
wire \ii2035|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5]|qx_net  ;
wire \ii2421|xy_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[12]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[21]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16]|qx_net  ;
wire \ii2796|xy_net  ;
wire \ii2806|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[25]_net  ;
wire \ii3282|xy_net  ;
wire \glue_dnum_s_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t85_out1_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[1]|qx_net  ;
wire \ii2737|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memwr_s_reg|qx_net  ;
wire \carry_12_ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[25]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3]|qx_net  ;
wire \ii2283|xy_net  ;
wire \ii2668|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[17]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5]|qx_net  ;
wire \ii2224|xy_net  ;
wire \carry_13_ADD_0|co_net  ;
wire \ii2599|xy_net  ;
wire \ii2609|xy_net  ;
wire \ii2610|xy_net  ;
wire \carry_9_4__ADD_0|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ;
wire \carry_9_7__ADD_3|co_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[22]|qx_net  ;
wire \carry_9_10__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4]|qx_net  ;
wire \ii2155|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]|qx_net  ;
wire \ii2926|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[6]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]|qx_net  ;
wire \ii2086|xy_net  ;
wire \ii2472|xy_net  ;
wire \ii2857|xy_net  ;
wire \ii3343|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14]|qx_net  ;
wire \ii2027|xy_net  ;
wire \ii2413|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16]|qx_net  ;
wire \ii2788|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59]|qx_net  ;
wire \carry_8_ADD_3|s_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1]|qx_net  ;
wire \ii2729|xy_net  ;
wire \ii2730|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[2]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10]|qx_net  ;
wire \carry_12_ADD_1|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17]|qx_net  ;
wire \ii2661|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net  ;
wire \carry_9_10__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[11]_net  ;
wire \ii2216|xy_net  ;
wire \ii2592|xy_net  ;
wire \ii2602|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26]|qx_net  ;
wire \carry_9_13__ADD_2|co_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[18]_net  ;
wire \ii2147|xy_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28]|qx_net  ;
wire \ii2918|xy_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf|xy_net  ;
wire \carry_9_11__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1]|qx_net  ;
wire \ii2078|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8]|qx_net  ;
wire \ii2464|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3]|qx_net  ;
wire \ii2849|xy_net  ;
wire \ii2850|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2]|qx_net  ;
wire \ii3335|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1]|qx_net  ;
wire \carry_8_ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_d_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[14]|qx_net  ;
wire \mipi_inst_u_mipi2|CM[7]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0]|qx_net  ;
wire \ii2781|xy_net  ;
wire \glue_rd_cmd_flag_reg|qx_net  ;
wire \carry_9_12__ADD_0|s_net  ;
wire \carry_12_ADD_5|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[9]_net  ;
wire \carry_9_5__ADD_7|co_net  ;
wire \ii2336|xy_net  ;
wire \ii2722|xy_net  ;
wire \carry_9_10__ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[18]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[4]_net  ;
wire \carry_12_1__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[8]_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf|xy_net  ;
wire \carry_9_13__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ;
wire \ii2653|xy_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[10]_net  ;
wire \glue_rx_packet_tx_packet_rstrf_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[2]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2]|qx_net  ;
wire \carry_9_11__ADD_4|s_net  ;
wire \ii2198|xy_net  ;
wire \ii2208|xy_net  ;
wire \ii2584|xy_net  ;
wire \u_8051_u_h6_8051|memdatao_comb[3]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[26]|qx_net  ;
wire \ii2139|xy_net  ;
wire \ii2140|xy_net  ;
wire \ii2525|xy_net  ;
wire \ii2911|xy_net  ;
wire \ii3386|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[7]_net  ;
wire \carry_9_12__ADD_4|s_net  ;
wire \carry_12_ADD_9|s_net  ;
wire \u_8051_u_h6_8051|memrd_comb_net  ;
wire \ii2071|xy_net  ;
wire \ii2456|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4]|qx_net  ;
wire \ii2842|xy_net  ;
wire \ii3327|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[25]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[15]_net  ;
wire \ii2773|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5]|qx_net  ;
wire \carry_9_13__ADD_4|s_net  ;
wire \u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17]|qx_net  ;
wire \carry_9_5__ADD_0|co_net  ;
wire \carry_9_8__ADD_3|co_net  ;
wire \ii2328|xy_net  ;
wire \ii2714|xy_net  ;
wire \carry_9_11__ADD_6|co_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[21]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13]|qx_net  ;
wire \glue_dnum_s_reg[12]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[8]_net  ;
wire \ii2645|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[6]_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg|qx_net  ;
wire \ii2191|xy_net  ;
wire \ii2201|xy_net  ;
wire \ii2576|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[9]|qx_net  ;
wire \ii2132|xy_net  ;
wire \ii2517|xy_net  ;
wire \ii2893|xy_net  ;
wire \ii2903|xy_net  ;
wire \ii3378|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[8]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4]|qx_net  ;
wire \ii2063|xy_net  ;
wire \ii2448|xy_net  ;
wire \ii2834|xy_net  ;
wire \ii3319|xy_net  ;
wire \ii3320|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[6]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25]|qx_net  ;
wire \glue_cmd_s_reg[3]|qx_net  ;
wire \ii2379|xy_net  ;
wire \ii2380|xy_net  ;
wire \ii2765|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[3]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2]|qx_net  ;
wire \ii2696|xy_net  ;
wire \ii2706|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3]|qx_net  ;
wire \glue_dnum_s_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[15]_net  ;
wire \mipi_inst_u_mipi2|prdata[19]_net  ;
wire \mipi_inst_u_mipi2|prdata[20]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1]|qx_net  ;
wire \ii2252|xy_net  ;
wire \ii2637|xy_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[19]_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[20]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[28]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3]|qx_net  ;
wire \ii2183|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6]|qx_net  ;
wire \ii2568|xy_net  ;
wire \carry_11_ADD_3|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[5]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[12]_net  ;
wire \ii2124|xy_net  ;
wire \ii2499|xy_net  ;
wire \ii2509|xy_net  ;
wire \ii2510|xy_net  ;
wire \ii2885|xy_net  ;
wire \ii3371|xy_net  ;
wire \carry_9_3__ADD_4|co_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[12]|qx_net  ;
wire \carry_9_6__ADD_7|co_net  ;
wire \ii2055|xy_net  ;
wire \glue_rd_cmd_flag_d_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7]|qx_net  ;
wire \ii2441|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18]|qx_net  ;
wire \ii2826|xy_net  ;
wire \ii3312|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_req_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[25]_net  ;
wire \carry_12_2__ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t86_out1_reg|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[1]_net  ;
wire \ii2372|xy_net  ;
wire \mcu_arbiter_u_emif2apb_memdatai_reg[3]|qx_net  ;
wire \ii2757|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net  ;
wire \carry_9_3__ADD_0|s_net  ;
wire \ii2688|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ;
wire \u_8051_u_h6_8051|port0o[1]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49]|qx_net  ;
wire \mipi_inst_u_mipi2|CO[1]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[14]_net  ;
wire \carry_11_ADD_7|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0]|qx_net  ;
wire \carry_8_ADD_6|co_net  ;
wire \ii2244|xy_net  ;
wire \ii2629|xy_net  ;
wire \ii2630|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net  ;
wire \carry_9_4__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[7]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6]|qx_net  ;
wire \ii2175|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6]|qx_net  ;
wire \ii2561|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7]|qx_net  ;
wire \carry_9_ADD_6|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30]|qx_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg|qx_net  ;
wire \ii2116|xy_net  ;
wire \ii2492|xy_net  ;
wire \ii2502|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0]|qx_net  ;
wire \ii2877|xy_net  ;
wire \ii3363|xy_net  ;
wire \carry_9_6__ADD_0|co_net  ;
wire \carry_9_5__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[7]_net  ;
wire \carry_9_9__ADD_3|co_net  ;
wire \carry_9_12__ADD_6|co_net  ;
wire \ii2047|xy_net  ;
wire \ii2433|xy_net  ;
wire \ii2818|xy_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[13]_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18]|qx_net  ;
wire \ii3304|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_rx_cmd[14]_net  ;
wire \carry_9_3__ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_write_data_temp_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[15]_net  ;
wire \glue_rx_packet_tx_packet_fifo_sync_readen_reg|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11]|qx_net  ;
wire \ii2749|xy_net  ;
wire \ii2750|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6]|qx_net  ;
wire \carry_9_6__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12]|qx_net  ;
wire \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19]|qx_net  ;
wire \ii2295|xy_net  ;
wire \ii2681|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7]|qx_net  ;
wire \ii3166|xy_net  ;
wire \mipi_inst_u_mipi2|CM[2]_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5]|qx_net  ;
wire \carry_9_4__ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_first_3e_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[4]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[5]_net  ;
wire \carry_9_7__ADD_0|s_net  ;
wire \ii2236|xy_net  ;
wire \ii2622|xy_net  ;
wire \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[13]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[3]_net  ;
wire \ii2167|xy_net  ;
wire \carry_9_5__ADD_4|s_net  ;
wire \mipi_inst_u_mipi2|prdata[6]_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3]|qx_net  ;
wire \carry_9_8__ADD_0|s_net  ;
wire \ii2108|xy_net  ;
wire \ii2098|xy_net  ;
wire \ii1998|xy_net  ;
wire \u_8051_u_h6_8051|memaddr_comb[4]_net  ;
wire \ii2484|xy_net  ;
wire \ii2870|xy_net  ;
wire \ii2869|xy_net  ;
wire \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[26]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3]|qx_net  ;
wire \mipi_inst_u_mipi1|periph_dphy_direction_net  ;
wire \ii3355|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4]|qx_net  ;
wire \carry_11_ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_rx_cmd_d_reg[3]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5]|qx_net  ;
wire \carry_9_6__ADD_4|s_net  ;
wire \ii2040|xy_net  ;
wire \ii2039|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[16]|qx_net  ;
wire \ii2425|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2]|qx_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[6]_net  ;
wire \ii2811|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ;
wire \carry_9_9__ADD_0|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[9]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[2]_net  ;
wire \ii2742|xy_net  ;
wire \carry_12_ADD_4|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7]|qx_net  ;
wire \carry_9_7__ADD_4|s_net  ;
wire \ii2287|xy_net  ;
wire \ii2673|xy_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[20]_net  ;
wire \mcu_arbiter_u_psram_u_psram|datao[19]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[10]_net  ;
wire \mcu_arbiter_code_sel_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4]|qx_net  ;
wire \carry_13_ADD_4|co_net  ;
wire \ii2228|xy_net  ;
wire \carry_9_4__ADD_4|co_net  ;
wire \ii2614|xy_net  ;
wire \carry_9_7__ADD_7|co_net  ;
wire \carry_9_8__ADD_4|s_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[11]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ;
wire \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7]|qx_net  ;
wire \carry_12_0__ADD_3|co_net  ;
wire \ii2160|xy_net  ;
wire \ii2159|xy_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[28]|qx_net  ;
wire \ii2931|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[10]_net  ;
wire \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[3]_net  ;
wire \ii1991|xy_net  ;
wire \ii2091|xy_net  ;
wire \ii2101|xy_net  ;
wire \carry_9_9__ADD_4|s_net  ;
wire \ii2476|xy_net  ;
wire \ii2862|xy_net  ;
wire \ii3347|xy_net  ;
wire \mcu_arbiter_reg_din_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7]|qx_net  ;
wire \carry_13_ADD_11|co_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[8]_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[0]|qx_net  ;
wire \ii2032|xy_net  ;
wire \ii2417|xy_net  ;
wire \ii2793|xy_net  ;
wire \ii2803|xy_net  ;
wire \carry_12_0__ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1]|qx_net  ;
wire \ii2734|xy_net  ;
wire \uut_dataReadBack_mipi_periph_tx_payload_reg[23]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15]|qx_net  ;
wire \mcu_arbiter_reg_memack_reg|qx_net  ;
wire \glue_dnum_s_reg[14]|qx_net  ;
wire \mipi_inst_u_mipi1|prdata[1]_net  ;
wire \carry_12_1__ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1]|qx_net  ;
wire \ii2665|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_rstsf_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10]|qx_net  ;
wire \ii2221|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ;
wire \ii2606|xy_net  ;
wire \ii2596|xy_net  ;
wire \carry_9_7__ADD_0|co_net  ;
wire \mcu_arbiter_func_reg[1]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3]|qx_net  ;
wire \carry_9_10__ADD_3|co_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[10]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4]|qx_net  ;
wire \carry_9_13__ADD_6|co_net  ;
wire \carry_12_2__ADD_4|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10]|qx_net  ;
wire \mipi_inst_u_mipi2|prdata[14]_net  ;
wire \ii2152|xy_net  ;
wire \ii2923|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[5]_net  ;
wire \carry_12_0__ADD_8|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12]|qx_net  ;
wire \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7]|qx_net  ;
wire \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[6]_net  ;
wire \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6]|qx_net  ;
wire \ii1983|xy_net  ;
wire \ii2083|xy_net  ;
wire \ii2468|xy_net  ;
wire \ii2854|xy_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[14]_net  ;
wire \mipi_inst_u_mipi1|periph_rx_payload[23]_net  ;
wire \ii3340|xy_net  ;
wire \ii3339|xy_net  ;
wire \mipi_inst_u_mipi2|prdata[27]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27]|qx_net  ;
wire \glue_cmd_s_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_rx_payload_d_reg[1]|qx_net  ;
wire \ii2410|xy_net  ;
wire \ii2409|xy_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_reg|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7]|qx_net  ;
wire \ii2785|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3]|qx_net  ;
wire \carry_12_1__ADD_8|s_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[27]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11]|qx_net  ;
wire \ii2341|xy_net  ;
wire \ii2726|xy_net  ;
wire \glue_dnum_s_reg[2]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[20]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[19]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3]|qx_net  ;
wire \ii2657|xy_net  ;
wire \carry_12_2__ADD_8|s_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4]|qx_net  ;
wire \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5]|qx_net  ;
wire \ii2213|xy_net  ;
wire \ii2588|xy_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0]|qx_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[11]_net  ;
wire \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40]|qx_net  ;
wire \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39]|qx_net  ;
wire \mcu_arbiter_u_pfifo_u_inst|dout[8]_net  ;
wire \ii2144|xy_net  ;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4] .always_en = 1;
LUT6 ii2686 (
	. xy ( \ii2686|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f1 ( \ii2685|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2686.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2686.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2686.config_data = 64'b0011000000000000001110100000000000110101000000000011111100000000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[6]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]|qx_net  ),
	. di ( \ii2480|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .PCK_LOCATION = "C16R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19]|qx_net  ),
	. di ( \ii2885|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .PLACE_LOCATION = "C6R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .PCK_LOCATION = "C6R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20]|qx_net  ),
	. di ( \ii2889|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .PLACE_LOCATION = "C8R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .PCK_LOCATION = "C8R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_13__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3] .always_en = 1;
LUT6 ii2687 (
	. xy ( \ii2687|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2612|xy_net  )
);
defparam ii2687.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2687.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2687.config_data = 64'b1110101011100000101010101010000001001010010000000000101000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .PCK_LOCATION = "C16R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3] .always_en = 1;
LUT6 ii2688 (
	. xy ( \ii2688|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \ii2612|xy_net  ),
	. f2 ( \ii2582|xy_net  ),
	. f1 ( \ii2687|xy_net  ),
	. f0 ( \ii2686|xy_net  )
);
defparam ii2688.PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.lut_0";
defparam ii2688.PCK_LOCATION = "C6R10.lp0.lut_0";
defparam ii2688.config_data = 64'b0101010101010101010001000100010101010101010101010100010001000100;
LUT6 ii2700 (
	. xy ( \ii2700|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2699|xy_net  )
);
defparam ii2700.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2700.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2700.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
LUT6 ii2690 (
	. xy ( \ii2690|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2689|xy_net  )
);
defparam ii2690.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2690.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2690.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
LUT6 ii2689 (
	. xy ( \ii2689|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2689.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2689.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2689.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[11]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[11] .always_en = 1;
LUT6 ii2701 (
	. xy ( \ii2701|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2701.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2701.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2701.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
LUT6 ii2691 (
	. xy ( \ii2691|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2691.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2691.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2691.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. di ( \ii2698|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[30]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[29]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2702 (
	. xy ( \ii2702|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]|qx_net  )
);
defparam ii2702.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2702.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2702.config_data = 64'b1011111110111100101100111011000010001111100011001000001110000000;
LUT6 ii2692 (
	. xy ( \ii2692|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]|qx_net  )
);
defparam ii2692.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2692.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2692.config_data = 64'b1011111110111100101100111011000010001111100011001000001110000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2] .always_en = 1;
LUT6 ii2703 (
	. xy ( \ii2703|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2702|xy_net  ),
	. f1 ( \ii2701|xy_net  ),
	. f0 ( \ii2700|xy_net  )
);
defparam ii2703.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2703.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2703.config_data = 64'b1111110011001100101010101010101011111100110011001010101010101010;
LUT6 ii2693 (
	. xy ( \ii2693|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2692|xy_net  ),
	. f1 ( \ii2691|xy_net  ),
	. f0 ( \ii2690|xy_net  )
);
defparam ii2693.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2693.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2693.config_data = 64'b1111110011001100101010101010101011111100110011001010101010101010;
LUT6 ii2704 (
	. xy ( \ii2704|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2704.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2704.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2704.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
LUT6 ii2694 (
	. xy ( \ii2694|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2694.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2694.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2694.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .PCK_LOCATION = "C10R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11] .always_en = 1;
LUT6 ii2705 (
	. xy ( \ii2705|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2705.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2705.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2705.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2695 (
	. xy ( \ii2695|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2695.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2695.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2695.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2706 (
	. xy ( \ii2706|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2705|xy_net  )
);
defparam ii2706.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2706.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2706.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
LUT6 ii2696 (
	. xy ( \ii2696|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2695|xy_net  )
);
defparam ii2696.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2696.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2696.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5] .always_en = 1;
LUT6 ii2707 (
	. xy ( \ii2707|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]|qx_net  )
);
defparam ii2707.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2707.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2707.config_data = 64'b1011111110111100101100111011000010001111100011001000001110000000;
LUT6 ii2697 (
	. xy ( \ii2697|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]|qx_net  )
);
defparam ii2697.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.lut_0";
defparam ii2697.PCK_LOCATION = "C8R8.lp0.lut_0";
defparam ii2697.config_data = 64'b1011111110111100101100111011000010001111100011001000001110000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_13__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21]|qx_net  ),
	. di ( \ii2891|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]|qx_net  ),
	. di ( \ii2481|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2] .always_en = 1;
LUT6 ii2708 (
	. xy ( \ii2708|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2707|xy_net  ),
	. f1 ( \ii2706|xy_net  ),
	. f0 ( \ii2704|xy_net  )
);
defparam ii2708.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2708.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2708.config_data = 64'b1111101010101010110011001100110011111010101010101100110011001100;
LUT6 ii2698 (
	. xy ( \ii2698|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2697|xy_net  ),
	. f1 ( \ii2696|xy_net  ),
	. f0 ( \ii2694|xy_net  )
);
defparam ii2698.PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.lut_0";
defparam ii2698.PCK_LOCATION = "C6R8.lp0.lut_0";
defparam ii2698.config_data = 64'b1111000010101010110011001100110011110000101010101100110011001100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .PCK_LOCATION = "C14R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .PCK_LOCATION = "C16R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[12]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[12] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27] .always_en = 1;
LUT6 ii2710 (
	. xy ( \ii2710|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]|qx_net  ),
	. f1 ( \ii2709|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2710.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.lut_0";
defparam ii2710.PCK_LOCATION = "C8R8.lp0.lut_0";
defparam ii2710.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
LUT6 ii2709 (
	. xy ( \ii2709|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2]|qx_net  )
);
defparam ii2709.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2709.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2709.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
LUT6 ii2699 (
	. xy ( \ii2699|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2699.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2699.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2699.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. di ( \ii2703|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28] .always_en = 1;
LUT6 ii2711 (
	. xy ( \ii2711|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2710|xy_net  )
);
defparam ii2711.PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.lut_0";
defparam ii2711.PCK_LOCATION = "C10R9.lp0.lut_0";
defparam ii2711.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
LUT6 u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly (
	. xy ( \u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly|xy_net  )
);
defparam u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp1.lut_0";
defparam u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly.PCK_LOCATION = "NONE";
defparam u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3] .always_en = 1;
LUT6 ii2712 (
	. xy ( \ii2712|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2712.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2712.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2712.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2713 (
	. xy ( \ii2713|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2712|xy_net  )
);
defparam ii2713.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2713.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2713.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .PCK_LOCATION = "C10R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4] .always_en = 1;
LUT6 ii2714 (
	. xy ( \ii2714|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2714.PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.lut_0";
defparam ii2714.PCK_LOCATION = "C6R10.lp0.lut_0";
defparam ii2714.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
LUT6 ii2715 (
	. xy ( \ii2715|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]|qx_net  )
);
defparam ii2715.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2715.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2715.config_data = 64'b1011111110111100101100111011000010001111100011001000001110000000;
LUT6 ii2716 (
	. xy ( \ii2716|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2715|xy_net  ),
	. f1 ( \ii2714|xy_net  ),
	. f0 ( \ii2713|xy_net  )
);
defparam ii2716.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2716.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2716.config_data = 64'b1111110011001100101010101010101011111100110011001010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]|qx_net  ),
	. di ( \ii2482|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22]|qx_net  ),
	. di ( \ii2893|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_13__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5] .always_en = 1;
LUT6 ii2717 (
	. xy ( \ii2717|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2717.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2717.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2717.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .PCK_LOCATION = "C16R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .PCK_LOCATION = "C14R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1] .always_en = 1;
LUT6 ii2718 (
	. xy ( \ii2718|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2717|xy_net  )
);
defparam ii2718.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2718.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2718.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[13]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[13] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_3__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0] .always_en = 1;
LUT6 ii2719 (
	. xy ( \ii2719|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2719.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.lut_0";
defparam ii2719.PCK_LOCATION = "C8R8.lp0.lut_0";
defparam ii2719.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
LUT6 ii2720 (
	. xy ( \ii2720|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]|qx_net  )
);
defparam ii2720.PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.lut_0";
defparam ii2720.PCK_LOCATION = "C10R9.lp0.lut_0";
defparam ii2720.config_data = 64'b1011111110111100101100111011000010001111100011001000001110000000;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10]|qx_net  ),
	. di ( \ii2585|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. di ( \ii2708|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. di ( \ii2716|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30] .always_en = 1;
LUT6 ii2721 (
	. xy ( \ii2721|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2720|xy_net  ),
	. f1 ( \ii2719|xy_net  ),
	. f0 ( \ii2718|xy_net  )
);
defparam ii2721.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2721.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2721.config_data = 64'b1111110011001100101010101010101011111100110011001010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4] .always_en = 1;
LUT6 ii2722 (
	. xy ( \ii2722|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2722.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam ii2722.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam ii2722.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2723 (
	. xy ( \ii2723|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \ii2722|xy_net  )
);
defparam ii2723.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2723.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2723.config_data = 64'b1111111110111011110000001000100000111111101110110000000010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .PLACE_LOCATION = "C14R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .PCK_LOCATION = "C14R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[0]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5] .always_en = 1;
LUT6 ii2724 (
	. xy ( \ii2724|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2724.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam ii2724.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam ii2724.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2725 (
	. xy ( \ii2725|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2725.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2725.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2725.config_data = 64'b1111011111100110110101011100010010110011101000101001000110000000;
LUT6 ii2726 (
	. xy ( \ii2726|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2725|xy_net  ),
	. f1 ( \ii2724|xy_net  ),
	. f0 ( \ii2723|xy_net  )
);
defparam ii2726.PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.lut_0";
defparam ii2726.PCK_LOCATION = "C6R10.lp0.lut_0";
defparam ii2726.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]|qx_net  ),
	. di ( \ii2483|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23]|qx_net  ),
	. di ( \ii2895|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_13__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6] .always_en = 1;
LUT6 ii2727 (
	. xy ( \ii2727|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2727.PLACE_LOCATION = "C4R12.le_tile.le_guts.lp0.lut_0";
defparam ii2727.PCK_LOCATION = "C4R12.lp0.lut_0";
defparam ii2727.config_data = 64'b1111111111110111111111011111010110001010100000101000100010000000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[19]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf.PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf.PCK_LOCATION = "C4R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[20]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .PCK_LOCATION = "C16R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .PCK_LOCATION = "C14R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2] .always_en = 1;
LUT6 ii2728 (
	. xy ( \ii2728|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f0 ( \ii2727|xy_net  )
);
defparam ii2728.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2728.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2728.config_data = 64'b0001000100010001000100010001000100110001000100010001000100010001;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[14]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[14] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_3__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1] .always_en = 1;
LUT6 ii2729 (
	. xy ( \ii2729|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2729.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2729.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2729.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2730 (
	. xy ( \ii2730|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2730.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2730.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2730.config_data = 64'b1111111001110110110111000101010010111010001100101001100000010000;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11]|qx_net  ),
	. di ( \ii2586|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. di ( \ii2721|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31] .always_en = 1;
LUT6 ii2731 (
	. xy ( \ii2731|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2730|xy_net  ),
	. f1 ( \ii2729|xy_net  ),
	. f0 ( \ii2728|xy_net  )
);
defparam ii2731.PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.lut_0";
defparam ii2731.PCK_LOCATION = "C6R10.lp0.lut_0";
defparam ii2731.config_data = 64'b0101000001000100010101010101010101010000010001000101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .PCK_LOCATION = "C8R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5] .always_en = 1;
LUT6 ii2732 (
	. xy ( \ii2732|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2732.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2732.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2732.config_data = 64'b1110111011001100001011100000110011100010110000000010001000000000;
LUT6 ii2733 (
	. xy ( \ii2733|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2733.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2733.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2733.config_data = 64'b1111101111101010011100110110001011011001110010000101000101000000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .PLACE_LOCATION = "C14R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .PCK_LOCATION = "C14R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[1]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6] .always_en = 1;
LUT6 ii2734 (
	. xy ( \ii2734|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f1 ( \ii2733|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2734.PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.lut_0";
defparam ii2734.PCK_LOCATION = "C6R10.lp0.lut_0";
defparam ii2734.config_data = 64'b1100111111000101110010101100000011001111110001011100101011000000;
LUT6 ii2735 (
	. xy ( \ii2735|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \ii2612|xy_net  ),
	. f2 ( \ii2582|xy_net  ),
	. f1 ( \ii2734|xy_net  ),
	. f0 ( \ii2732|xy_net  )
);
defparam ii2735.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2735.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2735.config_data = 64'b1100110011001100101010101010111111001100110011001010101010101010;
LUT6 ii2736 (
	. xy ( \ii2736|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2736.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2736.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2736.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]|qx_net  ),
	. di ( \ii2484|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24]|qx_net  ),
	. di ( \ii2897|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_13__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7] .always_en = 1;
LUT6 ii2737 (
	. xy ( \ii2737|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2737.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2737.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2737.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .PCK_LOCATION = "C16R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3] .always_en = 1;
LUT6 ii2738 (
	. xy ( \ii2738|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f2 ( \ii2737|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2738.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2738.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2738.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG glue_rx_packet_tx_packet_tx_hsync_fo_reg (
	. qx ( \glue_rx_packet_tx_packet_tx_hsync_fo_reg|qx_net  ),
	. di ( \ii2423|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.init = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_tx_hsync_fo_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[15]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[15] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_3__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2] .always_en = 1;
LUT6 ii2739 (
	. xy ( \ii2739|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2739.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2739.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2739.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
LUT6 ii2740 (
	. xy ( \ii2740|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2739|xy_net  ),
	. f1 ( \ii2738|xy_net  ),
	. f0 ( \ii2736|xy_net  )
);
defparam ii2740.PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.lut_0";
defparam ii2740.PCK_LOCATION = "C6R9.lp0.lut_0";
defparam ii2740.config_data = 64'b1111101010101010001100110011001111111010101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0]|qx_net  ),
	. di ( \ii2455|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12]|qx_net  ),
	. di ( \ii2587|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. di ( \ii2726|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32] .always_en = 1;
LUT6 ii2741 (
	. xy ( \ii2741|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2741.PLACE_LOCATION = "C4R10.le_tile.le_guts.lp0.lut_0";
defparam ii2741.PCK_LOCATION = "C4R10.lp0.lut_0";
defparam ii2741.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .PCK_LOCATION = "C8R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1] .always_en = 1;
LUT6 ii2742 (
	. xy ( \ii2742|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2742.PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.lut_0";
defparam ii2742.PCK_LOCATION = "C4R9.lp0.lut_0";
defparam ii2742.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
LUT6 ii2743 (
	. xy ( \ii2743|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f2 ( \ii2742|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2743.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2743.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2743.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .PLACE_LOCATION = "C14R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .PCK_LOCATION = "C14R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[2]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7] .always_en = 1;
LUT6 ii2744 (
	. xy ( \ii2744|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2744.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2744.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2744.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
LUT6 ii2745 (
	. xy ( \ii2745|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2744|xy_net  ),
	. f1 ( \ii2743|xy_net  ),
	. f0 ( \ii2741|xy_net  )
);
defparam ii2745.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.lut_0";
defparam ii2745.PCK_LOCATION = "C8R9.lp0.lut_0";
defparam ii2745.config_data = 64'b1111101010101010001100110011001111111010101010100011001100110011;
LUT6 ii2746 (
	. xy ( \ii2746|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2746.PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.lut_0";
defparam ii2746.PCK_LOCATION = "C6R10.lp0.lut_0";
defparam ii2746.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]|qx_net  ),
	. di ( \ii2485|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25]|qx_net  ),
	. di ( \ii2899|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net  ),
	. di ( \ii3021|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .PCK_LOCATION = "C16R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8] .always_en = 1;
LUT6 ii2747 (
	. xy ( \ii2747|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2747.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam ii2747.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam ii2747.config_data = 64'b1111010101110101100000000000000011110101011101011000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4] .always_en = 1;
LUT6 ii2748 (
	. xy ( \ii2748|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \ii2747|xy_net  ),
	. f0 ( \ii2612|xy_net  )
);
defparam ii2748.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2748.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2748.config_data = 64'b0001000100110001000100110011001100010001001100010001001100110011;
FIFO18K glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst (
	. dout ( {
		/* dout [63] (nc) */ nc0 ,
		/* dout [62] (nc) */ nc1 ,
		/* dout [61] (nc) */ nc2 ,
		/* dout [60] (nc) */ nc3 ,
		/* dout [59] (nc) */ nc4 ,
		/* dout [58] (nc) */ nc5 ,
		/* dout [57] (nc) */ nc6 ,
		/* dout [56] (nc) */ nc7 ,
		/* dout [55] (nc) */ nc8 ,
		/* dout [54] (nc) */ nc9 ,
		/* dout [53] (nc) */ nc10 ,
		/* dout [52] (nc) */ nc11 ,
		/* dout [51] (nc) */ nc12 ,
		/* dout [50] (nc) */ nc13 ,
		/* dout [49] (nc) */ nc14 ,
		/* dout [48] (nc) */ nc15 ,
		/* dout [47] (nc) */ nc16 ,
		/* dout [46] (nc) */ nc17 ,
		/* dout [45] (nc) */ nc18 ,
		/* dout [44] (nc) */ nc19 ,
		/* dout [43] (nc) */ nc20 ,
		/* dout [42] (nc) */ nc21 ,
		/* dout [41] (nc) */ nc22 ,
		/* dout [40] (nc) */ nc23 ,
		/* dout [39] (nc) */ nc24 ,
		/* dout [38] (nc) */ nc25 ,
		/* dout [37] (nc) */ nc26 ,
		/* dout [36] (nc) */ nc27 ,
		/* dout [35] (nc) */ nc28 ,
		/* dout [34] (nc) */ nc29 ,
		/* dout [33] (nc) */ nc30 ,
		/* dout [32] (nc) */ nc31 ,
		/* dout [31] (nc) */ nc32 ,
		/* dout [30] (nc) */ nc33 ,
		/* dout [29] (nc) */ nc34 ,
		/* dout [28] (nc) */ nc35 ,
		/* dout [27] (nc) */ nc36 ,
		/* dout [26] (nc) */ nc37 ,
		/* dout [25] (nc) */ nc38 ,
		/* dout [24] (nc) */ nc39 ,
		/* dout [23] (nc) */ nc40 ,
		/* dout [22] (nc) */ nc41 ,
		/* dout [21] (nc) */ nc42 ,
		/* dout [20] (nc) */ nc43 ,
		/* dout [19] (nc) */ nc44 ,
		/* dout [18] (nc) */ nc45 ,
		/* dout [17] (nc) */ nc46 ,
		/* dout [16] (nc) */ nc47 ,
		/* dout [15] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[15]_net ,
		/* dout [14] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[14]_net ,
		/* dout [13] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[13]_net ,
		/* dout [12] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[12]_net ,
		/* dout [11] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[11]_net ,
		/* dout [10] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[10]_net ,
		/* dout [9] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[9]_net ,
		/* dout [8] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[8]_net ,
		/* dout [7] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[7]_net ,
		/* dout [6] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[6]_net ,
		/* dout [5] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[5]_net ,
		/* dout [4] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[4]_net ,
		/* dout [3] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[3]_net ,
		/* dout [2] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[2]_net ,
		/* dout [1] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[1]_net ,
		/* dout [0] */ \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[0]_net 
	} ),
	. doutp ( )
,
	. din ( {
		/* din [63] */ \GND_0_inst|Y_net ,
		/* din [62] */ \GND_0_inst|Y_net ,
		/* din [61] */ \GND_0_inst|Y_net ,
		/* din [60] */ \GND_0_inst|Y_net ,
		/* din [59] */ \GND_0_inst|Y_net ,
		/* din [58] */ \GND_0_inst|Y_net ,
		/* din [57] */ \GND_0_inst|Y_net ,
		/* din [56] */ \GND_0_inst|Y_net ,
		/* din [55] */ \GND_0_inst|Y_net ,
		/* din [54] */ \GND_0_inst|Y_net ,
		/* din [53] */ \GND_0_inst|Y_net ,
		/* din [52] */ \GND_0_inst|Y_net ,
		/* din [51] */ \GND_0_inst|Y_net ,
		/* din [50] */ \GND_0_inst|Y_net ,
		/* din [49] */ \GND_0_inst|Y_net ,
		/* din [48] */ \GND_0_inst|Y_net ,
		/* din [47] */ \GND_0_inst|Y_net ,
		/* din [46] */ \GND_0_inst|Y_net ,
		/* din [45] */ \GND_0_inst|Y_net ,
		/* din [44] */ \GND_0_inst|Y_net ,
		/* din [43] */ \GND_0_inst|Y_net ,
		/* din [42] */ \GND_0_inst|Y_net ,
		/* din [41] */ \GND_0_inst|Y_net ,
		/* din [40] */ \GND_0_inst|Y_net ,
		/* din [39] */ \GND_0_inst|Y_net ,
		/* din [38] */ \GND_0_inst|Y_net ,
		/* din [37] */ \GND_0_inst|Y_net ,
		/* din [36] */ \GND_0_inst|Y_net ,
		/* din [35] */ \GND_0_inst|Y_net ,
		/* din [34] */ \GND_0_inst|Y_net ,
		/* din [33] */ \GND_0_inst|Y_net ,
		/* din [32] */ \GND_0_inst|Y_net ,
		/* din [31] */ \GND_0_inst|Y_net ,
		/* din [30] */ \GND_0_inst|Y_net ,
		/* din [29] */ \GND_0_inst|Y_net ,
		/* din [28] */ \GND_0_inst|Y_net ,
		/* din [27] */ \GND_0_inst|Y_net ,
		/* din [26] */ \GND_0_inst|Y_net ,
		/* din [25] */ \GND_0_inst|Y_net ,
		/* din [24] */ \GND_0_inst|Y_net ,
		/* din [23] */ \GND_0_inst|Y_net ,
		/* din [22] */ \GND_0_inst|Y_net ,
		/* din [21] */ \GND_0_inst|Y_net ,
		/* din [20] */ \GND_0_inst|Y_net ,
		/* din [19] */ \GND_0_inst|Y_net ,
		/* din [18] */ \GND_0_inst|Y_net ,
		/* din [17] */ \GND_0_inst|Y_net ,
		/* din [16] */ \GND_0_inst|Y_net ,
		/* din [15] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15]|qx_net ,
		/* din [14] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14]|qx_net ,
		/* din [13] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13]|qx_net ,
		/* din [12] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12]|qx_net ,
		/* din [11] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11]|qx_net ,
		/* din [10] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10]|qx_net ,
		/* din [9] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9]|qx_net ,
		/* din [8] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8]|qx_net ,
		/* din [7] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7]|qx_net ,
		/* din [6] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6]|qx_net ,
		/* din [5] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5]|qx_net ,
		/* din [4] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4]|qx_net ,
		/* din [3] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3]|qx_net ,
		/* din [2] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2]|qx_net ,
		/* din [1] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1]|qx_net ,
		/* din [0] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0]|qx_net 
	} ),
	. dinp ( {
		/* dinp [7] */ \GND_0_inst|Y_net ,
		/* dinp [6] */ \GND_0_inst|Y_net ,
		/* dinp [5] */ \GND_0_inst|Y_net ,
		/* dinp [4] */ \GND_0_inst|Y_net ,
		/* dinp [3] */ \GND_0_inst|Y_net ,
		/* dinp [2] */ \GND_0_inst|Y_net ,
		/* dinp [1] */ \GND_0_inst|Y_net ,
		/* dinp [0] */ \GND_0_inst|Y_net 
	} ),
	. writeclk ( \u_pll_pll_u0|CO0_net  ),
	. readclk ( \u_pll_pll_u0|CO0_net  ),
	. writeen ( \ii1990|xy_net  ),
	. readen ( \ii1989|xy_net  ),
	. reset ( \ii1987|xy_net  ),
	. regce ( \VCC_0_inst|Y_net  ),
	. writesave ( \GND_0_inst|Y_net  ),
	. writedrop ( \GND_0_inst|Y_net  ),
	. full ( ),
	. empty ( ),
	. almostfull ( ),
	. almostempty ( ),
	. overflow ( ),
	. underflow ( ),
	. eccoutdberr ( ),
	. eccoutsberr ( ),
	. eccreadaddr ( )
,
	. eccindberr ( \GND_0_inst|Y_net  ),
	. eccinsberr ( \GND_0_inst|Y_net  ),
	. writedropflag ( )
);
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.eccwriteen = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.writeclk_inv = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.eccreaden = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.readclk_inv = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.use_parity = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.outreg = 1;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.almostfullth = 988;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.almostemptyth = 512;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.writewidth = 18;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.readwidth = 18;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.peek = 1;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.PLACE_LOCATION = "C12R9.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst.PCK_LOCATION = "C12R9.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[16]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[16]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[16] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_3__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3] .always_en = 1;
LUT6 ii2749 (
	. xy ( \ii2749|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2749.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2749.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2749.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
LUT6 ii2750 (
	. xy ( \ii2750|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2749|xy_net  ),
	. f1 ( \ii2748|xy_net  ),
	. f0 ( \ii2746|xy_net  )
);
defparam ii2750.PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.lut_0";
defparam ii2750.PCK_LOCATION = "C8R10.lp0.lut_0";
defparam ii2750.config_data = 64'b1111101010101010001100110011001111111010101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1]|qx_net  ),
	. di ( \ii2456|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13]|qx_net  ),
	. di ( \ii2588|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. di ( \ii2731|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33] .always_en = 1;
LUT6 ii2751 (
	. xy ( \ii2751|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2751.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2751.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2751.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2] .always_en = 1;
LUT6 ii2752 (
	. xy ( \ii2752|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2752.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2752.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2752.config_data = 64'b1111010101110101100000000000000011110101011101011000000000000000;
LUT6 ii2753 (
	. xy ( \ii2753|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \ii2752|xy_net  ),
	. f0 ( \ii2612|xy_net  )
);
defparam ii2753.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2753.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2753.config_data = 64'b0001000100110001000100110011001100010001001100010001001100110011;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[10]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf.PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf.PCK_LOCATION = "C4R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[3]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[3] .always_en = 1;
LUT6 ii2754 (
	. xy ( \ii2754|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2754.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2754.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2754.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
LUT6 ii2755 (
	. xy ( \ii2755|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2754|xy_net  ),
	. f1 ( \ii2753|xy_net  ),
	. f0 ( \ii2751|xy_net  )
);
defparam ii2755.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2755.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2755.config_data = 64'b1111101010101010001100110011001111111010101010100011001100110011;
LUT6 ii2756 (
	. xy ( \ii2756|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2756.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2756.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2756.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]|qx_net  ),
	. di ( \ii2486|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26]|qx_net  ),
	. di ( \ii2901|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .PLACE_LOCATION = "C6R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .PCK_LOCATION = "C6R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0] .always_en = 1;
LUT6 ii2757 (
	. xy ( \ii2757|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2757.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2757.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2757.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5] .always_en = 1;
LUT6 ii2758 (
	. xy ( \ii2758|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f2 ( \ii2757|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2758.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2758.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2758.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG mcu_arbiter_fifo_clr_d_reg (
	. qx ( \mcu_arbiter_fifo_clr_d_reg|qx_net  ),
	. di ( \mcu_arbiter_fifo_clr_s_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_fifo_clr_d_reg.latch_mode = 0;
defparam mcu_arbiter_fifo_clr_d_reg.init = 0;
defparam mcu_arbiter_fifo_clr_d_reg.PLACE_LOCATION = "C4R23.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_fifo_clr_d_reg.sr_inv = 1;
defparam mcu_arbiter_fifo_clr_d_reg.sync_mode = 0;
defparam mcu_arbiter_fifo_clr_d_reg.no_sr = 0;
defparam mcu_arbiter_fifo_clr_d_reg.sr_value = 0;
defparam mcu_arbiter_fifo_clr_d_reg.PCK_LOCATION = "C4R23.lp0.reg0";
defparam mcu_arbiter_fifo_clr_d_reg.clk_inv = 0;
defparam mcu_arbiter_fifo_clr_d_reg.en_inv = 0;
defparam mcu_arbiter_fifo_clr_d_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[17]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[17]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[17] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_3__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4] .always_en = 1;
LUT6 ii2759 (
	. xy ( \ii2759|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2759.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2759.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2759.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
LUT6 ii2760 (
	. xy ( \ii2760|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2759|xy_net  ),
	. f1 ( \ii2758|xy_net  ),
	. f0 ( \ii2756|xy_net  )
);
defparam ii2760.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2760.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2760.config_data = 64'b1111101010101010001100110011001111111010101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2]|qx_net  ),
	. di ( \ii2457|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14]|qx_net  ),
	. di ( \ii2589|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. di ( \ii2735|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34] .always_en = 1;
LUT6 ii2761 (
	. xy ( \ii2761|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3]|qx_net  )
);
defparam ii2761.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2761.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2761.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3] .always_en = 1;
LUT6 ii2762 (
	. xy ( \ii2762|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]|qx_net  ),
	. f1 ( \ii2761|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2762.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2762.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2762.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
LUT6 ii2763 (
	. xy ( \ii2763|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2762|xy_net  )
);
defparam ii2763.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2763.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2763.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[4]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[4] .always_en = 1;
LUT6 ii2764 (
	. xy ( \ii2764|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2764.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2764.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2764.config_data = 64'b1000101000001010100000100000001010001000000010001000000000000000;
LUT6 ii2765 (
	. xy ( \ii2765|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f2 ( \ii2764|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2765.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2765.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2765.config_data = 64'b0000111000001111000011100000111100001110000011110000111000001111;
REG glue_rd_cmd_flag_d_reg (
	. qx ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. di ( \glue_rd_cmd_flag_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rd_cmd_flag_d_reg.latch_mode = 0;
defparam glue_rd_cmd_flag_d_reg.init = 0;
defparam glue_rd_cmd_flag_d_reg.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam glue_rd_cmd_flag_d_reg.sr_inv = 1;
defparam glue_rd_cmd_flag_d_reg.sync_mode = 0;
defparam glue_rd_cmd_flag_d_reg.no_sr = 0;
defparam glue_rd_cmd_flag_d_reg.sr_value = 0;
defparam glue_rd_cmd_flag_d_reg.PCK_LOCATION = "C14R27.lp0.reg0";
defparam glue_rd_cmd_flag_d_reg.clk_inv = 0;
defparam glue_rd_cmd_flag_d_reg.en_inv = 0;
defparam glue_rd_cmd_flag_d_reg.always_en = 1;
LUT6 ii2766 (
	. xy ( \ii2766|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2766.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2766.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2766.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
LUT6 ii2767 (
	. xy ( \ii2767|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2767.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2767.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2767.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27]|qx_net  ),
	. di ( \ii2903|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .PLACE_LOCATION = "C8R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .PCK_LOCATION = "C8R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2] .always_en = 1;
LUT6 ii2768 (
	. xy ( \ii2768|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2767|xy_net  ),
	. f1 ( \ii2766|xy_net  ),
	. f0 ( \ii2765|xy_net  )
);
defparam ii2768.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2768.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2768.config_data = 64'b1111110011001100010101010101010111111100110011000101010101010101;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6] .always_en = 1;
LUT6 ii2770 (
	. xy ( \ii2770|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2770.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam ii2770.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam ii2770.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
LUT6 ii2769 (
	. xy ( \ii2769|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2769.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam ii2769.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam ii2769.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_3__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[18]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[18]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[18] .always_en = 1;
LUT6 ii2771 (
	. xy ( \ii2771|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f2 ( \ii2770|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2771.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2771.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2771.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. di ( \ii2740|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15]|qx_net  ),
	. di ( \ii2590|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3]|qx_net  ),
	. di ( \ii2458|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[3] .always_en = 1;
LUT6 ii2772 (
	. xy ( \ii2772|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2772.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2772.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2772.config_data = 64'b1111101111101010110110011100100001110011011000100101000101000000;
LUT6 ii2773 (
	. xy ( \ii2773|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2772|xy_net  ),
	. f1 ( \ii2771|xy_net  ),
	. f0 ( \ii2769|xy_net  )
);
defparam ii2773.PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.lut_0";
defparam ii2773.PCK_LOCATION = "C8R11.lp0.lut_0";
defparam ii2773.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2774 (
	. xy ( \ii2774|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2774.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2774.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2774.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc48 ,
		/* a_mac_out [23] (nc) */ nc49 ,
		/* a_mac_out [22] (nc) */ nc50 ,
		/* a_mac_out [21] (nc) */ nc51 ,
		/* a_mac_out [20] (nc) */ nc52 ,
		/* a_mac_out [19] (nc) */ nc53 ,
		/* a_mac_out [18] (nc) */ nc54 ,
		/* a_mac_out [17] (nc) */ nc55 ,
		/* a_mac_out [16] (nc) */ nc56 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc57 ,
		/* a_mac_out [2] (nc) */ nc58 ,
		/* a_mac_out [1] (nc) */ nc59 ,
		/* a_mac_out [0] (nc) */ nc60 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.PLACE_LOCATION = "C22R19.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.PCK_LOCATION = "C22R19.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[5]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18] .always_en = 1;
REG mcu_arbiter_code_sel_reg (
	. qx ( \mcu_arbiter_code_sel_reg|qx_net  ),
	. di ( \ii3318|xy_net  ),
	. sr ( ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_code_sel_reg.latch_mode = 0;
defparam mcu_arbiter_code_sel_reg.init = 0;
defparam mcu_arbiter_code_sel_reg.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_code_sel_reg.sr_inv = 0;
defparam mcu_arbiter_code_sel_reg.sync_mode = 1;
defparam mcu_arbiter_code_sel_reg.no_sr = 1;
defparam mcu_arbiter_code_sel_reg.sr_value = 0;
defparam mcu_arbiter_code_sel_reg.PCK_LOCATION = "C4R18.lp0.reg0";
defparam mcu_arbiter_code_sel_reg.clk_inv = 0;
defparam mcu_arbiter_code_sel_reg.en_inv = 0;
defparam mcu_arbiter_code_sel_reg.always_en = 1;
LUT6 ii2775 (
	. xy ( \ii2775|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2775.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam ii2775.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam ii2775.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
LUT6 ii2776 (
	. xy ( \ii2776|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f2 ( \ii2775|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2776.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2776.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2776.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
LUT6 ii2777 (
	. xy ( \ii2777|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2777.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2777.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2777.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28]|qx_net  ),
	. di ( \ii2905|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3] .always_en = 1;
REG glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.PCK_LOCATION = "C4R6.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg.always_en = 1;
LUT6 ii2778 (
	. xy ( \ii2778|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2777|xy_net  ),
	. f1 ( \ii2776|xy_net  ),
	. f0 ( \ii2774|xy_net  )
);
defparam ii2778.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2778.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2778.config_data = 64'b1111000001010101001100110011001111110000010101010011001100110011;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7] .always_en = 1;
REG mcu_arbiter_mipi_sel_reg (
	. qx ( \mcu_arbiter_mipi_sel_reg|qx_net  ),
	. di ( \ii3322|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_mipi_sel_reg.latch_mode = 0;
defparam mcu_arbiter_mipi_sel_reg.init = 0;
defparam mcu_arbiter_mipi_sel_reg.PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_mipi_sel_reg.sr_inv = 1;
defparam mcu_arbiter_mipi_sel_reg.sync_mode = 0;
defparam mcu_arbiter_mipi_sel_reg.no_sr = 0;
defparam mcu_arbiter_mipi_sel_reg.sr_value = 0;
defparam mcu_arbiter_mipi_sel_reg.PCK_LOCATION = "C4R14.lp0.reg0";
defparam mcu_arbiter_mipi_sel_reg.clk_inv = 0;
defparam mcu_arbiter_mipi_sel_reg.en_inv = 0;
defparam mcu_arbiter_mipi_sel_reg.always_en = 1;
LUT6 ii2780 (
	. xy ( \ii2780|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2780.PLACE_LOCATION = "C4R12.le_tile.le_guts.lp0.lut_0";
defparam ii2780.PCK_LOCATION = "C4R12.lp0.lut_0";
defparam ii2780.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2779 (
	. xy ( \ii2779|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2779.PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.lut_0";
defparam ii2779.PCK_LOCATION = "C4R13.lp0.lut_0";
defparam ii2779.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_3__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[19]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[19]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[20]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[20]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[20] .always_en = 1;
LUT6 ii2781 (
	. xy ( \ii2781|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f2 ( \ii2780|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2781.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2781.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2781.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. di ( \ii2745|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16]|qx_net  ),
	. di ( \ii2591|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4]|qx_net  ),
	. di ( \ii2459|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4] .always_en = 1;
LUT6 ii2782 (
	. xy ( \ii2782|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2782.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2782.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2782.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2783 (
	. xy ( \ii2783|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2782|xy_net  ),
	. f1 ( \ii2781|xy_net  ),
	. f0 ( \ii2779|xy_net  )
);
defparam ii2783.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2783.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2783.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2784 (
	. xy ( \ii2784|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2784.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2784.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2784.config_data = 64'b0011000100100000001100010010000000110001001000000011000100100000;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[6]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20] .always_en = 1;
LUT6 ii2785 (
	. xy ( \ii2785|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2785.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii2785.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii2785.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2786 (
	. xy ( \ii2786|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f2 ( \ii2785|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2786.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam ii2786.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam ii2786.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
LUT6 ii2787 (
	. xy ( \ii2787|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2787.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2787.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2787.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30]|qx_net  ),
	. di ( \ii2911|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29]|qx_net  ),
	. di ( \ii2907|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4] .always_en = 1;
LUT6 ii2788 (
	. xy ( \ii2788|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2787|xy_net  ),
	. f1 ( \ii2786|xy_net  ),
	. f0 ( \ii2784|xy_net  )
);
defparam ii2788.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2788.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2788.config_data = 64'b1111101010101010001100110011001111111010101010100011001100110011;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8] .always_en = 1;
LUT6 ii2800 (
	. xy ( \ii2800|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2800.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2800.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2800.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2790 (
	. xy ( \ii2790|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2790.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam ii2790.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam ii2790.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2789 (
	. xy ( \ii2789|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2789.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam ii2789.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam ii2789.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_3__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .PLACE_LOCATION = "C6R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .PCK_LOCATION = "C6R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[21]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[21]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[21] .always_en = 1;
LUT6 ii2801 (
	. xy ( \ii2801|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f2 ( \ii2800|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2801.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2801.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2801.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
LUT6 ii2791 (
	. xy ( \ii2791|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f2 ( \ii2790|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2791.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2791.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2791.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. di ( \ii2750|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17]|qx_net  ),
	. di ( \ii2592|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5]|qx_net  ),
	. di ( \ii2460|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5] .always_en = 1;
LUT6 ii2802 (
	. xy ( \ii2802|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2802.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2802.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2802.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2792 (
	. xy ( \ii2792|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2792.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2792.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2792.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2803 (
	. xy ( \ii2803|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2802|xy_net  ),
	. f1 ( \ii2801|xy_net  ),
	. f0 ( \ii2799|xy_net  )
);
defparam ii2803.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.lut_0";
defparam ii2803.PCK_LOCATION = "C18R12.lp0.lut_0";
defparam ii2803.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2793 (
	. xy ( \ii2793|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2792|xy_net  ),
	. f1 ( \ii2791|xy_net  ),
	. f0 ( \ii2789|xy_net  )
);
defparam ii2793.PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.lut_0";
defparam ii2793.PCK_LOCATION = "C8R12.lp0.lut_0";
defparam ii2793.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2804 (
	. xy ( \ii2804|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2804.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam ii2804.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam ii2804.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
LUT6 ii2794 (
	. xy ( \ii2794|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2794.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2794.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2794.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .PCK_LOCATION = "C16R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[7]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[7] .always_en = 1;
REG glue_rx_packet_tx_packet_sc1_rstf_reg (
	. qx ( \glue_rx_packet_tx_packet_sc1_rstf_reg|qx_net  ),
	. di ( \ii2422|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.init = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.PCK_LOCATION = "C20R7.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_sc1_rstf_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21] .always_en = 1;
LUT6 ii2805 (
	. xy ( \ii2805|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2805.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2805.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2805.config_data = 64'b1000000010001000100000101000101011110101111111011111011111111111;
LUT6 ii2795 (
	. xy ( \ii2795|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2795.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam ii2795.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam ii2795.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2806 (
	. xy ( \ii2806|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f2 ( \ii2805|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2806.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.lut_0";
defparam ii2806.PCK_LOCATION = "C18R12.lp0.lut_0";
defparam ii2806.config_data = 64'b1101000011110000110100001111000011010000111100001101000011110000;
LUT6 ii2796 (
	. xy ( \ii2796|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f2 ( \ii2795|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2796.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2796.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2796.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
ADD1_A carry_9_4__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_4__ADD_0|co_net  ),
	. s ( \carry_9_4__ADD_0|s_net  )
);
defparam carry_9_4__ADD_0.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_0.a_inv = "true";
defparam carry_9_4__ADD_0.PCK_LOCATION = "C8R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0] .always_en = 1;
LUT6 ii2807 (
	. xy ( \ii2807|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2807.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2807.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2807.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2797 (
	. xy ( \ii2797|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2797.PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.lut_0";
defparam ii2797.PCK_LOCATION = "C14R11.lp0.lut_0";
defparam ii2797.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31]|qx_net  ),
	. di ( \ii2913|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5] .always_en = 1;
ADD1_A carry_9_4__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1]|qx_net  ),
	. ci ( \carry_9_4__ADD_0|co_net  ),
	. co ( \carry_9_4__ADD_1|co_net  ),
	. s ( \carry_9_4__ADD_1|s_net  )
);
defparam carry_9_4__ADD_1.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_1.a_inv = "true";
defparam carry_9_4__ADD_1.PCK_LOCATION = "C8R8.lp0.add2.add0";
LUT6 ii2808 (
	. xy ( \ii2808|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2807|xy_net  ),
	. f1 ( \ii2806|xy_net  ),
	. f0 ( \ii2804|xy_net  )
);
defparam ii2808.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2808.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2808.config_data = 64'b1111000001010101001100110011001111110000010101010011001100110011;
LUT6 ii2798 (
	. xy ( \ii2798|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2797|xy_net  ),
	. f1 ( \ii2796|xy_net  ),
	. f0 ( \ii2794|xy_net  )
);
defparam ii2798.PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.lut_0";
defparam ii2798.PCK_LOCATION = "C14R12.lp0.lut_0";
defparam ii2798.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
ADD1_A carry_9_4__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2]|qx_net  ),
	. ci ( \carry_9_4__ADD_1|co_net  ),
	. co ( \carry_9_4__ADD_2|co_net  ),
	. s ( \carry_9_4__ADD_2|s_net  )
);
defparam carry_9_4__ADD_2.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_2.a_inv = "true";
defparam carry_9_4__ADD_2.PCK_LOCATION = "C8R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9] .always_en = 1;
REG \mcu_arbiter_func_reg[0]  (
	. qx ( \mcu_arbiter_func_reg[0]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[0] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[0] .init = 0;
defparam \mcu_arbiter_func_reg[0] .PLACE_LOCATION = "C8R17.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[0] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[0] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[0] .no_sr = 0;
defparam \mcu_arbiter_func_reg[0] .sr_value = 0;
defparam \mcu_arbiter_func_reg[0] .PCK_LOCATION = "C8R17.lp0.reg0";
defparam \mcu_arbiter_func_reg[0] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[0] .en_inv = 0;
defparam \mcu_arbiter_func_reg[0] .always_en = 0;
LUT6 ii2810 (
	. xy ( \ii2810|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2810.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam ii2810.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam ii2810.config_data = 64'b0000101000000010000010000000000000001010000000100000100000000000;
LUT6 ii2809 (
	. xy ( \ii2809|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2809.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2809.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2809.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2799 (
	. xy ( \ii2799|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2799.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2799.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2799.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net  ),
	. di ( \ii3050|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8] .always_en = 1;
ADD1_A carry_9_4__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3]|qx_net  ),
	. ci ( \carry_9_4__ADD_2|co_net  ),
	. co ( \carry_9_4__ADD_3|co_net  ),
	. s ( \carry_9_4__ADD_3|s_net  )
);
defparam carry_9_4__ADD_3.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_3.a_inv = "true";
defparam carry_9_4__ADD_3.PCK_LOCATION = "C8R8.lp0.add2.add0";
GND GND_0_inst (
	. Y ( \GND_0_inst|Y_net  )
);
defparam GND_0_inst.PLACE_LOCATION = "NONE";
defparam GND_0_inst.PCK_LOCATION = "NONE";
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[22]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[22]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[22] .always_en = 1;
LUT6 ii2811 (
	. xy ( \ii2811|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f2 ( \ii2810|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2811.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2811.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2811.config_data = 64'b0000110000001110000011010000111100001100000011100000110100001111;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. di ( \ii2755|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18]|qx_net  ),
	. di ( \ii2593|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18] .always_en = 1;
ADD1_A carry_9_4__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4]|qx_net  ),
	. ci ( \carry_9_4__ADD_3|co_net  ),
	. co ( \carry_9_4__ADD_4|co_net  ),
	. s ( \carry_9_4__ADD_4|s_net  )
);
defparam carry_9_4__ADD_4.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_4.a_inv = "true";
defparam carry_9_4__ADD_4.PCK_LOCATION = "C8R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6]|qx_net  ),
	. di ( \ii2461|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6] .always_en = 1;
LUT6 ii2812 (
	. xy ( \ii2812|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2812.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.lut_0";
defparam ii2812.PCK_LOCATION = "C10R12.lp0.lut_0";
defparam ii2812.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc61 ,
		/* a_mac_out [23] (nc) */ nc62 ,
		/* a_mac_out [22] (nc) */ nc63 ,
		/* a_mac_out [21] (nc) */ nc64 ,
		/* a_mac_out [20] (nc) */ nc65 ,
		/* a_mac_out [19] (nc) */ nc66 ,
		/* a_mac_out [18] (nc) */ nc67 ,
		/* a_mac_out [17] (nc) */ nc68 ,
		/* a_mac_out [16] (nc) */ nc69 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc70 ,
		/* a_mac_out [2] (nc) */ nc71 ,
		/* a_mac_out [1] (nc) */ nc72 ,
		/* a_mac_out [0] (nc) */ nc73 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.PLACE_LOCATION = "C22R21.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.PCK_LOCATION = "C22R21.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0.amac_output_mode = 0;
ADD1_A carry_9_4__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5]|qx_net  ),
	. ci ( \carry_9_4__ADD_4|co_net  ),
	. co ( \carry_9_4__ADD_5|co_net  ),
	. s ( \carry_9_4__ADD_5|s_net  )
);
defparam carry_9_4__ADD_5.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_5.a_inv = "true";
defparam carry_9_4__ADD_5.PCK_LOCATION = "C8R8.lp0.add2.add0";
REG glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg|qx_net  ),
	. di ( \ii2427|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.PCK_LOCATION = "C16R10.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg.always_en = 1;
LUT6 ii2813 (
	. xy ( \ii2813|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2812|xy_net  ),
	. f1 ( \ii2811|xy_net  ),
	. f0 ( \ii2809|xy_net  )
);
defparam ii2813.PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.lut_0";
defparam ii2813.PCK_LOCATION = "C10R11.lp0.lut_0";
defparam ii2813.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
ADD1_A carry_9_4__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6]|qx_net  ),
	. ci ( \carry_9_4__ADD_5|co_net  ),
	. co ( \carry_9_4__ADD_6|co_net  ),
	. s ( \carry_9_4__ADD_6|s_net  )
);
defparam carry_9_4__ADD_6.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_6.a_inv = "true";
defparam carry_9_4__ADD_6.PCK_LOCATION = "C8R8.lp0.add2.add0";
VCC VCC_0_inst (
	. Y ( \VCC_0_inst|Y_net  )
);
defparam VCC_0_inst.PLACE_LOCATION = "NONE";
defparam VCC_0_inst.PCK_LOCATION = "NONE";
LUT6 ii2814 (
	. xy ( \ii2814|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4]|qx_net  )
);
defparam ii2814.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2814.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2814.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1] .always_en = 1;
ADD1_A carry_9_4__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7]|qx_net  ),
	. ci ( \carry_9_4__ADD_6|co_net  ),
	. co ( \carry_9_4__ADD_7|co_net  ),
	. s ( \carry_9_4__ADD_7|s_net  )
);
defparam carry_9_4__ADD_7.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_7.a_inv = "true";
defparam carry_9_4__ADD_7.PCK_LOCATION = "C8R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[8]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22] .always_en = 1;
LUT6 ii2815 (
	. xy ( \ii2815|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]|qx_net  ),
	. f1 ( \ii2814|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2815.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2815.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2815.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
ADD1_A carry_9_4__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_4__ADD_7|co_net  ),
	. co ( \carry_9_4__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_4__ADD_8.PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_4__ADD_8.a_inv = "false";
defparam carry_9_4__ADD_8.PCK_LOCATION = "C8R9.lp0.add2.add0";
LUT6 ii2816 (
	. xy ( \ii2816|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[4]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2815|xy_net  )
);
defparam ii2816.PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.lut_0";
defparam ii2816.PCK_LOCATION = "C14R10.lp0.lut_0";
defparam ii2816.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1] .always_en = 1;
LUT6 ii2817 (
	. xy ( \ii2817|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2817.PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.lut_0";
defparam ii2817.PCK_LOCATION = "C14R13.lp0.lut_0";
defparam ii2817.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6] .always_en = 1;
LUT6 ii2818 (
	. xy ( \ii2818|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2818.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2818.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2818.config_data = 64'b1000000010001000100000101000101011110101111111011111011111111111;
REG \mcu_arbiter_func_reg[1]  (
	. qx ( \mcu_arbiter_func_reg[1]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[1] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[1] .init = 0;
defparam \mcu_arbiter_func_reg[1] .PLACE_LOCATION = "C4R17.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[1] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[1] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[1] .no_sr = 0;
defparam \mcu_arbiter_func_reg[1] .sr_value = 0;
defparam \mcu_arbiter_func_reg[1] .PCK_LOCATION = "C4R17.lp0.reg0";
defparam \mcu_arbiter_func_reg[1] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[1] .en_inv = 0;
defparam \mcu_arbiter_func_reg[1] .always_en = 0;
LUT6 ii2820 (
	. xy ( \ii2820|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2820.PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.lut_0";
defparam ii2820.PCK_LOCATION = "C14R12.lp0.lut_0";
defparam ii2820.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2819 (
	. xy ( \ii2819|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f2 ( \ii2818|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2819.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2819.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2819.config_data = 64'b1101000011110000110100001111000011010000111100001101000011110000;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[23]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[23]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[23] .always_en = 1;
LUT6 ii2821 (
	. xy ( \ii2821|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2820|xy_net  ),
	. f1 ( \ii2819|xy_net  ),
	. f0 ( \ii2817|xy_net  )
);
defparam ii2821.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2821.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2821.config_data = 64'b1111000001010101001100110011001111110000010101010011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. di ( \ii2768|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. di ( \ii2760|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20]|qx_net  ),
	. di ( \ii2596|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .PLACE_LOCATION = "C10R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .PCK_LOCATION = "C10R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19]|qx_net  ),
	. di ( \ii2594|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .PLACE_LOCATION = "C10R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .PCK_LOCATION = "C10R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7]|qx_net  ),
	. di ( \ii2462|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7] .always_en = 1;
LUT6 ii2822 (
	. xy ( \ii2822|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2822.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam ii2822.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam ii2822.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2823 (
	. xy ( \ii2823|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2823.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam ii2823.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam ii2823.config_data = 64'b0000101000000010000010000000000000001010000000100000100000000000;
REG glue_rx_packet_tx_packet_u_scaler_t50_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.PLACE_LOCATION = "C20R26.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.PCK_LOCATION = "C20R26.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t50_out1_reg.always_en = 1;
LUT6 ii2824 (
	. xy ( \ii2824|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f2 ( \ii2823|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2824.PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.lut_0";
defparam ii2824.PCK_LOCATION = "C14R12.lp0.lut_0";
defparam ii2824.config_data = 64'b0000110000001110000011010000111100001100000011100000110100001111;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[9]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23] .always_en = 1;
LUT6 ii2825 (
	. xy ( \ii2825|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2825.PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.lut_0";
defparam ii2825.PCK_LOCATION = "C14R12.lp0.lut_0";
defparam ii2825.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2826 (
	. xy ( \ii2826|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2825|xy_net  ),
	. f1 ( \ii2824|xy_net  ),
	. f0 ( \ii2822|xy_net  )
);
defparam ii2826.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2826.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2826.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.PCK_LOCATION = "C20R15.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg.always_en = 1;
LUT6 ii2827 (
	. xy ( \ii2827|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2827.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2827.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2827.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7] .always_en = 1;
LUT6 ii2828 (
	. xy ( \ii2828|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2828.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam ii2828.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam ii2828.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \mcu_arbiter_func_reg[2]  (
	. qx ( \mcu_arbiter_func_reg[2]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[2] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[2] .init = 0;
defparam \mcu_arbiter_func_reg[2] .PLACE_LOCATION = "C4R17.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[2] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[2] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[2] .no_sr = 0;
defparam \mcu_arbiter_func_reg[2] .sr_value = 0;
defparam \mcu_arbiter_func_reg[2] .PCK_LOCATION = "C4R17.lp0.reg0";
defparam \mcu_arbiter_func_reg[2] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[2] .en_inv = 0;
defparam \mcu_arbiter_func_reg[2] .always_en = 0;
LUT6 ii2830 (
	. xy ( \ii2830|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2830.PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.lut_0";
defparam ii2830.PCK_LOCATION = "C14R12.lp0.lut_0";
defparam ii2830.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2829 (
	. xy ( \ii2829|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f2 ( \ii2828|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2829.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2829.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2829.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[24]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[24]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[24] .always_en = 1;
LUT6 ii2831 (
	. xy ( \ii2831|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2830|xy_net  ),
	. f1 ( \ii2829|xy_net  ),
	. f0 ( \ii2827|xy_net  )
);
defparam ii2831.PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.lut_0";
defparam ii2831.PCK_LOCATION = "C14R13.lp0.lut_0";
defparam ii2831.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. di ( \ii2773|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21]|qx_net  ),
	. di ( \ii2597|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .PLACE_LOCATION = "C10R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .PCK_LOCATION = "C10R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21] .always_en = 1;
LUT6 ii2832 (
	. xy ( \ii2832|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2832.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2832.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2832.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2833 (
	. xy ( \ii2833|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2833.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2833.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2833.config_data = 64'b0000101000000010000010000000000000001010000000100000100000000000;
REG glue_rx_packet_tx_packet_rx_cmd_valid_d_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_valid_d_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd_valid_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.PCK_LOCATION = "C4R8.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_d_reg.always_en = 1;
LUT6 ii2834 (
	. xy ( \ii2834|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f2 ( \ii2833|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2834.PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.lut_0";
defparam ii2834.PCK_LOCATION = "C14R13.lp0.lut_0";
defparam ii2834.config_data = 64'b0000110000001110000011010000111100001100000011100000110100001111;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .PCK_LOCATION = "C16R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24] .always_en = 1;
LUT6 ii2835 (
	. xy ( \ii2835|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2835.PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.lut_0";
defparam ii2835.PCK_LOCATION = "C14R12.lp0.lut_0";
defparam ii2835.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
ADD1_A carry_13_ADD_10 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10]|qx_net  ),
	. ci ( \carry_13_ADD_9|co_net  ),
	. co ( \carry_13_ADD_10|co_net  ),
	. s ( \carry_13_ADD_10|s_net  )
);
defparam carry_13_ADD_10.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_10.a_inv = "false";
defparam carry_13_ADD_10.PCK_LOCATION = "C18R22.lp0.add2.add0";
LUT6 ii2836 (
	. xy ( \ii2836|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2835|xy_net  ),
	. f1 ( \ii2834|xy_net  ),
	. f0 ( \ii2832|xy_net  )
);
defparam ii2836.PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.lut_0";
defparam ii2836.PCK_LOCATION = "C14R13.lp0.lut_0";
defparam ii2836.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
ADD1_A carry_13_ADD_11 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]|qx_net  ),
	. ci ( \carry_13_ADD_10|co_net  ),
	. co ( \carry_13_ADD_11|co_net  ),
	. s ( \carry_13_ADD_11|s_net  )
);
defparam carry_13_ADD_11.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_11.a_inv = "false";
defparam carry_13_ADD_11.PCK_LOCATION = "C18R22.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3] .always_en = 1;
LUT6 ii2837 (
	. xy ( \ii2837|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2837.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam ii2837.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam ii2837.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8] .always_en = 1;
ADD1_A carry_13_ADD_12 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \GND_0_inst|Y_net  ),
	. ci ( \carry_13_ADD_11|co_net  ),
	. co ( ),
	. s ( \carry_13_ADD_12|s_net  )
);
defparam carry_13_ADD_12.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_12.a_inv = "false";
defparam carry_13_ADD_12.PCK_LOCATION = "C18R22.lp0.add2.add0";
LUT6 ii2838 (
	. xy ( \ii2838|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2838.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam ii2838.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam ii2838.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \mcu_arbiter_func_reg[3]  (
	. qx ( \mcu_arbiter_func_reg[3]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[3] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[3] .init = 0;
defparam \mcu_arbiter_func_reg[3] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[3] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[3] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[3] .no_sr = 0;
defparam \mcu_arbiter_func_reg[3] .sr_value = 0;
defparam \mcu_arbiter_func_reg[3] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_func_reg[3] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[3] .en_inv = 0;
defparam \mcu_arbiter_func_reg[3] .always_en = 0;
LUT6 ii2840 (
	. xy ( \ii2840|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2840.PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.lut_0";
defparam ii2840.PCK_LOCATION = "C14R13.lp0.lut_0";
defparam ii2840.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
LUT6 ii2839 (
	. xy ( \ii2839|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f2 ( \ii2838|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2839.PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.lut_0";
defparam ii2839.PCK_LOCATION = "C14R14.lp0.lut_0";
defparam ii2839.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[25]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[25]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[25] .always_en = 1;
LUT6 ii2841 (
	. xy ( \ii2841|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2840|xy_net  ),
	. f1 ( \ii2839|xy_net  ),
	. f0 ( \ii2837|xy_net  )
);
defparam ii2841.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam ii2841.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam ii2841.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. di ( \ii2778|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22]|qx_net  ),
	. di ( \ii2598|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .PLACE_LOCATION = "C10R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .PCK_LOCATION = "C10R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22] .always_en = 1;
LUT6 ii2842 (
	. xy ( \ii2842|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2842.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2842.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2842.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_8__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0] .always_en = 1;
LUT6 ii2843 (
	. xy ( \ii2843|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2843.PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.lut_0";
defparam ii2843.PCK_LOCATION = "C8R13.lp0.lut_0";
defparam ii2843.config_data = 64'b0000101000000010000010000000000000001010000000100000100000000000;
REG glue_rx_packet_tx_packet_sc1_fifo_readen_reg (
	. qx ( \glue_rx_packet_tx_packet_sc1_fifo_readen_reg|qx_net  ),
	. di ( \ii2339|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.init = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.PCK_LOCATION = "C16R9.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_sc1_fifo_readen_reg.always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[2]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf.PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf.PCK_LOCATION = "C4R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2844 (
	. xy ( \ii2844|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f2 ( \ii2843|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2844.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2844.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2844.config_data = 64'b0000110000001110000011010000111100001100000011100000110100001111;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .PCK_LOCATION = "C16R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25] .always_en = 1;
LUT6 ii2845 (
	. xy ( \ii2845|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2845.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2845.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2845.config_data = 64'b1111011110110011111001101010001011010101100100011100010010000000;
REG glue_rx_packet_tx_packet_rx_active_hs_d_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_active_hs_d_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|RxActiveHS_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.PCK_LOCATION = "C4R6.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_active_hs_d_reg.always_en = 1;
SIO io_phone_rst_inst (
	. f_id ( {
		/* f_id [1] (nc) */ nc74 ,
		/* f_id [0] */ \io_phone_rst_inst|f_id[0]_net 
	} ),
	. clk_en ( ),
	. fclk ( ),
	. od ( )
,
	. oen ( ),
	. rstn ( ),
	. setn ( ),
	. PAD ( phone_rst )
);
defparam io_phone_rst_inst.DDR_PREG_EN = 0;
defparam io_phone_rst_inst.FCLK_GATE_EN = 0;
defparam io_phone_rst_inst.FOEN_SEL = 0;
defparam io_phone_rst_inst.RSTN_SYNC = 0;
defparam io_phone_rst_inst.OUT_SEL = 0;
defparam io_phone_rst_inst.DDR_EN = 0;
defparam io_phone_rst_inst.NDR = 0;
defparam io_phone_rst_inst.VPCI_EN = 0;
defparam io_phone_rst_inst.ID_RSTN_EN = 0;
defparam io_phone_rst_inst.KEEP = 0;
defparam io_phone_rst_inst.PDR = 0;
defparam io_phone_rst_inst.SETN_INV = 0;
defparam io_phone_rst_inst.SETN_SYNC = 0;
defparam io_phone_rst_inst.FIN_SEL = 0;
defparam io_phone_rst_inst.ID_SETN_EN = 0;
defparam io_phone_rst_inst.DDR_REG_EN = 0;
defparam io_phone_rst_inst.FOUT_SEL = 0;
defparam io_phone_rst_inst.OEN_RSTN_EN = 0;
defparam io_phone_rst_inst.NS_LV = 3;
defparam io_phone_rst_inst.optional_function = "";
defparam io_phone_rst_inst.OD_RSTN_EN = 0;
defparam io_phone_rst_inst.RSTN_INV = 0;
defparam io_phone_rst_inst.is_clk_io = "false";
defparam io_phone_rst_inst.PLACE_LOCATION = "C24R11.io_guts.iob_ck.I0.I60.Iioc1";
defparam io_phone_rst_inst.OEN_SETN_EN = 0;
defparam io_phone_rst_inst.OEN_SEL = 0;
defparam io_phone_rst_inst.PCK_LOCATION = "NONE";
defparam io_phone_rst_inst.OD_SETN_EN = 0;
defparam io_phone_rst_inst.CLK_INV = 0;
defparam io_phone_rst_inst.is_signal_monitor_io = 1'b0;
defparam io_phone_rst_inst.DDR_NREG_EN = 0;
defparam io_phone_rst_inst.RX_DIG_EN = 1;
LUT6 ii2846 (
	. xy ( \ii2846|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2845|xy_net  ),
	. f1 ( \ii2844|xy_net  ),
	. f0 ( \ii2842|xy_net  )
);
defparam ii2846.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii2846.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii2846.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4] .always_en = 1;
LUT6 ii2847 (
	. xy ( \ii2847|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5]|qx_net  )
);
defparam ii2847.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2847.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2847.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0]|qx_net  ),
	. di ( \ii2471|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .PCK_LOCATION = "C6R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[0] .always_en = 1;
LUT6 ii2848 (
	. xy ( \ii2848|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]|qx_net  ),
	. f1 ( \ii2847|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2848.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2848.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2848.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[25]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \mcu_arbiter_func_reg[4]  (
	. qx ( \mcu_arbiter_func_reg[4]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[4] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[4] .init = 0;
defparam \mcu_arbiter_func_reg[4] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[4] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[4] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[4] .no_sr = 0;
defparam \mcu_arbiter_func_reg[4] .sr_value = 0;
defparam \mcu_arbiter_func_reg[4] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_func_reg[4] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[4] .en_inv = 0;
defparam \mcu_arbiter_func_reg[4] .always_en = 0;
LUT6 ii2850 (
	. xy ( \ii2850|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6]|qx_net  )
);
defparam ii2850.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2850.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2850.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
LUT6 ii2849 (
	. xy ( \ii2849|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[5]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2848|xy_net  )
);
defparam ii2849.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2849.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2849.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[26]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[26]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[26] .always_en = 1;
LUT6 ii2851 (
	. xy ( \ii2851|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]|qx_net  ),
	. f1 ( \ii2850|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2851.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2851.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2851.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. di ( \ii2783|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .PCK_LOCATION = "C6R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23]|qx_net  ),
	. di ( \ii2599|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .PLACE_LOCATION = "C10R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .PCK_LOCATION = "C10R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23] .always_en = 1;
LUT6 ii2852 (
	. xy ( \ii2852|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[6]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2851|xy_net  )
);
defparam ii2852.PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.lut_0";
defparam ii2852.PCK_LOCATION = "C14R11.lp0.lut_0";
defparam ii2852.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_8__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1] .always_en = 1;
LUT6 ii2853 (
	. xy ( \ii2853|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7]|qx_net  )
);
defparam ii2853.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2853.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2853.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
EMB18K glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0 (
	. doa ( {
		/* doa [63] (nc) */ nc75 ,
		/* doa [62] (nc) */ nc76 ,
		/* doa [61] (nc) */ nc77 ,
		/* doa [60] (nc) */ nc78 ,
		/* doa [59] (nc) */ nc79 ,
		/* doa [58] (nc) */ nc80 ,
		/* doa [57] (nc) */ nc81 ,
		/* doa [56] (nc) */ nc82 ,
		/* doa [55] (nc) */ nc83 ,
		/* doa [54] (nc) */ nc84 ,
		/* doa [53] (nc) */ nc85 ,
		/* doa [52] (nc) */ nc86 ,
		/* doa [51] (nc) */ nc87 ,
		/* doa [50] (nc) */ nc88 ,
		/* doa [49] (nc) */ nc89 ,
		/* doa [48] (nc) */ nc90 ,
		/* doa [47] (nc) */ nc91 ,
		/* doa [46] (nc) */ nc92 ,
		/* doa [45] (nc) */ nc93 ,
		/* doa [44] (nc) */ nc94 ,
		/* doa [43] (nc) */ nc95 ,
		/* doa [42] (nc) */ nc96 ,
		/* doa [41] (nc) */ nc97 ,
		/* doa [40] (nc) */ nc98 ,
		/* doa [39] (nc) */ nc99 ,
		/* doa [38] (nc) */ nc100 ,
		/* doa [37] (nc) */ nc101 ,
		/* doa [36] (nc) */ nc102 ,
		/* doa [35] (nc) */ nc103 ,
		/* doa [34] (nc) */ nc104 ,
		/* doa [33] (nc) */ nc105 ,
		/* doa [32] (nc) */ nc106 ,
		/* doa [31] (nc) */ nc107 ,
		/* doa [30] (nc) */ nc108 ,
		/* doa [29] (nc) */ nc109 ,
		/* doa [28] (nc) */ nc110 ,
		/* doa [27] (nc) */ nc111 ,
		/* doa [26] (nc) */ nc112 ,
		/* doa [25] (nc) */ nc113 ,
		/* doa [24] (nc) */ nc114 ,
		/* doa [23] (nc) */ nc115 ,
		/* doa [22] (nc) */ nc116 ,
		/* doa [21] (nc) */ nc117 ,
		/* doa [20] (nc) */ nc118 ,
		/* doa [19] (nc) */ nc119 ,
		/* doa [18] (nc) */ nc120 ,
		/* doa [17] (nc) */ nc121 ,
		/* doa [16] (nc) */ nc122 ,
		/* doa [15] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[15]_net ,
		/* doa [14] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[14]_net ,
		/* doa [13] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[13]_net ,
		/* doa [12] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[12]_net ,
		/* doa [11] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[11]_net ,
		/* doa [10] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[10]_net ,
		/* doa [9] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[9]_net ,
		/* doa [8] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[8]_net ,
		/* doa [7] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[7]_net ,
		/* doa [6] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[6]_net ,
		/* doa [5] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[5]_net ,
		/* doa [4] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[4]_net ,
		/* doa [3] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[3]_net ,
		/* doa [2] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[2]_net ,
		/* doa [1] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[1]_net ,
		/* doa [0] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[0]_net 
	} ),
	. dob ( )
,
	. dopa ( )
,
	. dopb ( )
,
	. addra ( {
		/* addra [13] */ \GND_0_inst|Y_net ,
		/* addra [12] */ \GND_0_inst|Y_net ,
		/* addra [11] */ \GND_0_inst|Y_net ,
		/* addra [10] */ \GND_0_inst|Y_net ,
		/* addra [9] */ \ii2035|xy_net ,
		/* addra [8] */ \ii2034|xy_net ,
		/* addra [7] */ \ii2033|xy_net ,
		/* addra [6] */ \ii2032|xy_net ,
		/* addra [5] */ \ii2031|xy_net ,
		/* addra [4] */ \ii2030|xy_net ,
		/* addra [3] */ \ii2029|xy_net ,
		/* addra [2] */ \ii2028|xy_net ,
		/* addra [1] */ \ii2027|xy_net ,
		/* addra [0] */ \ii2026|xy_net 
	} ),
	. addrb ( {
		/* addrb [13] */ \GND_0_inst|Y_net ,
		/* addrb [12] */ \GND_0_inst|Y_net ,
		/* addrb [11] */ \GND_0_inst|Y_net ,
		/* addrb [10] */ \GND_0_inst|Y_net ,
		/* addrb [9] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9]|qx_net ,
		/* addrb [8] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8]|qx_net ,
		/* addrb [7] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7]|qx_net ,
		/* addrb [6] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6]|qx_net ,
		/* addrb [5] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5]|qx_net ,
		/* addrb [4] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4]|qx_net ,
		/* addrb [3] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3]|qx_net ,
		/* addrb [2] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2]|qx_net ,
		/* addrb [1] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1]|qx_net ,
		/* addrb [0] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0]|qx_net 
	} ),
	. clka ( \u_pll_pll_u0|CO0_net  ),
	. clkb ( \u_pll_pll_u0|CO0_net  ),
	. dia ( )
,
	. dib ( {
		/* dib [63] (nc) */ nc123 ,
		/* dib [62] (nc) */ nc124 ,
		/* dib [61] (nc) */ nc125 ,
		/* dib [60] (nc) */ nc126 ,
		/* dib [59] (nc) */ nc127 ,
		/* dib [58] (nc) */ nc128 ,
		/* dib [57] (nc) */ nc129 ,
		/* dib [56] (nc) */ nc130 ,
		/* dib [55] (nc) */ nc131 ,
		/* dib [54] (nc) */ nc132 ,
		/* dib [53] (nc) */ nc133 ,
		/* dib [52] (nc) */ nc134 ,
		/* dib [51] (nc) */ nc135 ,
		/* dib [50] (nc) */ nc136 ,
		/* dib [49] (nc) */ nc137 ,
		/* dib [48] (nc) */ nc138 ,
		/* dib [47] (nc) */ nc139 ,
		/* dib [46] (nc) */ nc140 ,
		/* dib [45] (nc) */ nc141 ,
		/* dib [44] (nc) */ nc142 ,
		/* dib [43] (nc) */ nc143 ,
		/* dib [42] (nc) */ nc144 ,
		/* dib [41] (nc) */ nc145 ,
		/* dib [40] (nc) */ nc146 ,
		/* dib [39] (nc) */ nc147 ,
		/* dib [38] (nc) */ nc148 ,
		/* dib [37] (nc) */ nc149 ,
		/* dib [36] (nc) */ nc150 ,
		/* dib [35] (nc) */ nc151 ,
		/* dib [34] (nc) */ nc152 ,
		/* dib [33] (nc) */ nc153 ,
		/* dib [32] (nc) */ nc154 ,
		/* dib [31] (nc) */ nc155 ,
		/* dib [30] (nc) */ nc156 ,
		/* dib [29] (nc) */ nc157 ,
		/* dib [28] (nc) */ nc158 ,
		/* dib [27] (nc) */ nc159 ,
		/* dib [26] (nc) */ nc160 ,
		/* dib [25] (nc) */ nc161 ,
		/* dib [24] (nc) */ nc162 ,
		/* dib [23] (nc) */ nc163 ,
		/* dib [22] (nc) */ nc164 ,
		/* dib [21] (nc) */ nc165 ,
		/* dib [20] (nc) */ nc166 ,
		/* dib [19] (nc) */ nc167 ,
		/* dib [18] (nc) */ nc168 ,
		/* dib [17] (nc) */ nc169 ,
		/* dib [16] (nc) */ nc170 ,
		/* dib [15] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15]|qx_net ,
		/* dib [14] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14]|qx_net ,
		/* dib [13] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13]|qx_net ,
		/* dib [12] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12]|qx_net ,
		/* dib [11] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11]|qx_net ,
		/* dib [10] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10]|qx_net ,
		/* dib [9] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9]|qx_net ,
		/* dib [8] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8]|qx_net ,
		/* dib [7] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7]|qx_net ,
		/* dib [6] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6]|qx_net ,
		/* dib [5] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5]|qx_net ,
		/* dib [4] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4]|qx_net ,
		/* dib [3] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3]|qx_net ,
		/* dib [2] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2]|qx_net ,
		/* dib [1] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1]|qx_net ,
		/* dib [0] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0]|qx_net 
	} ),
	. dipa ( )
,
	. dipb ( )
,
	. cea ( \VCC_0_inst|Y_net  ),
	. ceb ( \VCC_0_inst|Y_net  ),
	. regcea ( \VCC_0_inst|Y_net  ),
	. regceb ( ),
	. regsra ( \VCC_0_inst|Y_net  ),
	. regsrb ( ),
	. wea ( {
		/* wea [3] */ \GND_0_inst|Y_net ,
		/* wea [2] */ \GND_0_inst|Y_net ,
		/* wea [1] */ \GND_0_inst|Y_net ,
		/* wea [0] */ \GND_0_inst|Y_net 
	} ),
	. web ( {
		/* web [3] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net ,
		/* web [2] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net ,
		/* web [1] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net ,
		/* web [0] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net 
	} ),
	. eccoutdberr ( ),
	. eccoutsberr ( ),
	. eccreadaddr ( )
,
	. eccindberr ( \GND_0_inst|Y_net  ),
	. eccinsberr ( \GND_0_inst|Y_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_1d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_1e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_1f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.eccreaden = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_00 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_01 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_02 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_2a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.emb5k_1_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_03 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_2b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_04 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_2c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_05 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_2d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_06 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_2e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_07 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_2f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_08 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_09 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_10 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_11 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.PCK_LOCATION = "C12R13.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.outreg_a = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_12 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_3a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.outreg_b = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_13 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_3b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.clkb_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_14 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_3c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.eccwriteen = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_15 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_3d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_16 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_00 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_3e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_17 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_01 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_3f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_18 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_02 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_20 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.rammode = "sdp";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.use_parity = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_19 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_03 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_21 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_04 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_22 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.emb5k_2_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_05 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_23 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_06 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_24 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.initp_07 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_25 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_26 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_27 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_28 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_30 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_29 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_31 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_32 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_33 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_34 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_35 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_36 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_37 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_38 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_39 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.emb5k_3_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.extension_mode = "power";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.clka_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.width_a = 18;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.writemode_a = "write_first";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.width_b = 18;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.writemode_b = "write_first";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_0a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_0b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_0c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_0d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_0e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.emb5k_4_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_0f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.PLACE_LOCATION = "C12R13.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_1a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_1b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0.init_1c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
LUT6 ii2854 (
	. xy ( \ii2854|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]|qx_net  ),
	. f1 ( \ii2853|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2854.PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.lut_0";
defparam ii2854.PCK_LOCATION = "C14R10.lp0.lut_0";
defparam ii2854.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
EMB18K glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1 (
	. doa ( {
		/* doa [63] (nc) */ nc171 ,
		/* doa [62] (nc) */ nc172 ,
		/* doa [61] (nc) */ nc173 ,
		/* doa [60] (nc) */ nc174 ,
		/* doa [59] (nc) */ nc175 ,
		/* doa [58] (nc) */ nc176 ,
		/* doa [57] (nc) */ nc177 ,
		/* doa [56] (nc) */ nc178 ,
		/* doa [55] (nc) */ nc179 ,
		/* doa [54] (nc) */ nc180 ,
		/* doa [53] (nc) */ nc181 ,
		/* doa [52] (nc) */ nc182 ,
		/* doa [51] (nc) */ nc183 ,
		/* doa [50] (nc) */ nc184 ,
		/* doa [49] (nc) */ nc185 ,
		/* doa [48] (nc) */ nc186 ,
		/* doa [47] (nc) */ nc187 ,
		/* doa [46] (nc) */ nc188 ,
		/* doa [45] (nc) */ nc189 ,
		/* doa [44] (nc) */ nc190 ,
		/* doa [43] (nc) */ nc191 ,
		/* doa [42] (nc) */ nc192 ,
		/* doa [41] (nc) */ nc193 ,
		/* doa [40] (nc) */ nc194 ,
		/* doa [39] (nc) */ nc195 ,
		/* doa [38] (nc) */ nc196 ,
		/* doa [37] (nc) */ nc197 ,
		/* doa [36] (nc) */ nc198 ,
		/* doa [35] (nc) */ nc199 ,
		/* doa [34] (nc) */ nc200 ,
		/* doa [33] (nc) */ nc201 ,
		/* doa [32] (nc) */ nc202 ,
		/* doa [31] (nc) */ nc203 ,
		/* doa [30] (nc) */ nc204 ,
		/* doa [29] (nc) */ nc205 ,
		/* doa [28] (nc) */ nc206 ,
		/* doa [27] (nc) */ nc207 ,
		/* doa [26] (nc) */ nc208 ,
		/* doa [25] (nc) */ nc209 ,
		/* doa [24] (nc) */ nc210 ,
		/* doa [23] (nc) */ nc211 ,
		/* doa [22] (nc) */ nc212 ,
		/* doa [21] (nc) */ nc213 ,
		/* doa [20] (nc) */ nc214 ,
		/* doa [19] (nc) */ nc215 ,
		/* doa [18] (nc) */ nc216 ,
		/* doa [17] (nc) */ nc217 ,
		/* doa [16] (nc) */ nc218 ,
		/* doa [15] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[15]_net ,
		/* doa [14] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[14]_net ,
		/* doa [13] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[13]_net ,
		/* doa [12] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[12]_net ,
		/* doa [11] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[11]_net ,
		/* doa [10] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[10]_net ,
		/* doa [9] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[9]_net ,
		/* doa [8] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[8]_net ,
		/* doa [7] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[7]_net ,
		/* doa [6] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[6]_net ,
		/* doa [5] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[5]_net ,
		/* doa [4] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[4]_net ,
		/* doa [3] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[3]_net ,
		/* doa [2] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[2]_net ,
		/* doa [1] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[1]_net ,
		/* doa [0] */ \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[0]_net 
	} ),
	. dob ( )
,
	. dopa ( )
,
	. dopb ( )
,
	. addra ( {
		/* addra [13] */ \GND_0_inst|Y_net ,
		/* addra [12] */ \GND_0_inst|Y_net ,
		/* addra [11] */ \GND_0_inst|Y_net ,
		/* addra [10] */ \GND_0_inst|Y_net ,
		/* addra [9] */ \ii2035|xy_net ,
		/* addra [8] */ \ii2034|xy_net ,
		/* addra [7] */ \ii2033|xy_net ,
		/* addra [6] */ \ii2032|xy_net ,
		/* addra [5] */ \ii2031|xy_net ,
		/* addra [4] */ \ii2030|xy_net ,
		/* addra [3] */ \ii2029|xy_net ,
		/* addra [2] */ \ii2028|xy_net ,
		/* addra [1] */ \ii2027|xy_net ,
		/* addra [0] */ \ii2026|xy_net 
	} ),
	. addrb ( {
		/* addrb [13] */ \GND_0_inst|Y_net ,
		/* addrb [12] */ \GND_0_inst|Y_net ,
		/* addrb [11] */ \GND_0_inst|Y_net ,
		/* addrb [10] */ \GND_0_inst|Y_net ,
		/* addrb [9] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9]|qx_net ,
		/* addrb [8] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8]|qx_net ,
		/* addrb [7] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7]|qx_net ,
		/* addrb [6] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6]|qx_net ,
		/* addrb [5] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5]|qx_net ,
		/* addrb [4] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4]|qx_net ,
		/* addrb [3] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3]|qx_net ,
		/* addrb [2] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2]|qx_net ,
		/* addrb [1] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1]|qx_net ,
		/* addrb [0] */ \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0]|qx_net 
	} ),
	. clka ( \u_pll_pll_u0|CO0_net  ),
	. clkb ( \u_pll_pll_u0|CO0_net  ),
	. dia ( )
,
	. dib ( {
		/* dib [63] (nc) */ nc219 ,
		/* dib [62] (nc) */ nc220 ,
		/* dib [61] (nc) */ nc221 ,
		/* dib [60] (nc) */ nc222 ,
		/* dib [59] (nc) */ nc223 ,
		/* dib [58] (nc) */ nc224 ,
		/* dib [57] (nc) */ nc225 ,
		/* dib [56] (nc) */ nc226 ,
		/* dib [55] (nc) */ nc227 ,
		/* dib [54] (nc) */ nc228 ,
		/* dib [53] (nc) */ nc229 ,
		/* dib [52] (nc) */ nc230 ,
		/* dib [51] (nc) */ nc231 ,
		/* dib [50] (nc) */ nc232 ,
		/* dib [49] (nc) */ nc233 ,
		/* dib [48] (nc) */ nc234 ,
		/* dib [47] (nc) */ nc235 ,
		/* dib [46] (nc) */ nc236 ,
		/* dib [45] (nc) */ nc237 ,
		/* dib [44] (nc) */ nc238 ,
		/* dib [43] (nc) */ nc239 ,
		/* dib [42] (nc) */ nc240 ,
		/* dib [41] (nc) */ nc241 ,
		/* dib [40] (nc) */ nc242 ,
		/* dib [39] (nc) */ nc243 ,
		/* dib [38] (nc) */ nc244 ,
		/* dib [37] (nc) */ nc245 ,
		/* dib [36] (nc) */ nc246 ,
		/* dib [35] (nc) */ nc247 ,
		/* dib [34] (nc) */ nc248 ,
		/* dib [33] (nc) */ nc249 ,
		/* dib [32] (nc) */ nc250 ,
		/* dib [31] (nc) */ nc251 ,
		/* dib [30] (nc) */ nc252 ,
		/* dib [29] (nc) */ nc253 ,
		/* dib [28] (nc) */ nc254 ,
		/* dib [27] (nc) */ nc255 ,
		/* dib [26] (nc) */ nc256 ,
		/* dib [25] (nc) */ nc257 ,
		/* dib [24] (nc) */ nc258 ,
		/* dib [23] (nc) */ nc259 ,
		/* dib [22] (nc) */ nc260 ,
		/* dib [21] (nc) */ nc261 ,
		/* dib [20] (nc) */ nc262 ,
		/* dib [19] (nc) */ nc263 ,
		/* dib [18] (nc) */ nc264 ,
		/* dib [17] (nc) */ nc265 ,
		/* dib [16] (nc) */ nc266 ,
		/* dib [15] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31]|qx_net ,
		/* dib [14] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30]|qx_net ,
		/* dib [13] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29]|qx_net ,
		/* dib [12] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28]|qx_net ,
		/* dib [11] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27]|qx_net ,
		/* dib [10] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26]|qx_net ,
		/* dib [9] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25]|qx_net ,
		/* dib [8] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24]|qx_net ,
		/* dib [7] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23]|qx_net ,
		/* dib [6] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22]|qx_net ,
		/* dib [5] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21]|qx_net ,
		/* dib [4] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20]|qx_net ,
		/* dib [3] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19]|qx_net ,
		/* dib [2] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18]|qx_net ,
		/* dib [1] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17]|qx_net ,
		/* dib [0] */ \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16]|qx_net 
	} ),
	. dipa ( )
,
	. dipb ( )
,
	. cea ( \VCC_0_inst|Y_net  ),
	. ceb ( \VCC_0_inst|Y_net  ),
	. regcea ( \VCC_0_inst|Y_net  ),
	. regceb ( ),
	. regsra ( \VCC_0_inst|Y_net  ),
	. regsrb ( ),
	. wea ( {
		/* wea [3] */ \GND_0_inst|Y_net ,
		/* wea [2] */ \GND_0_inst|Y_net ,
		/* wea [1] */ \GND_0_inst|Y_net ,
		/* wea [0] */ \GND_0_inst|Y_net 
	} ),
	. web ( {
		/* web [3] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net ,
		/* web [2] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net ,
		/* web [1] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net ,
		/* web [0] */ \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net 
	} ),
	. eccoutdberr ( ),
	. eccoutsberr ( ),
	. eccreadaddr ( )
,
	. eccindberr ( \GND_0_inst|Y_net  ),
	. eccinsberr ( \GND_0_inst|Y_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_1d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_1e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_1f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.eccreaden = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_00 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_01 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_02 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_2a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.emb5k_1_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_03 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_2b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_04 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_2c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_05 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_2d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_06 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_2e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_07 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_2f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_08 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_09 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_10 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_11 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.PCK_LOCATION = "C12R17.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.outreg_a = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_12 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_3a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.outreg_b = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_13 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_3b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.clkb_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_14 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_3c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.eccwriteen = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_15 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_3d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_16 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_00 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_3e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_17 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_01 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_3f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_18 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_02 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_20 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.rammode = "sdp";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.use_parity = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_19 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_03 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_21 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_04 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_22 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.emb5k_2_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_05 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_23 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_06 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_24 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.initp_07 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_25 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_26 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_27 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_28 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_30 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_29 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_31 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_32 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_33 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_34 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_35 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_36 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_37 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_38 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_39 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.emb5k_3_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.extension_mode = "power";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.clka_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.width_a = 18;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.writemode_a = "write_first";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.width_b = 18;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.writemode_b = "write_first";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_0a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_0b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_0c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_0d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_0e = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.emb5k_4_init_file = "none";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_0f = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.PLACE_LOCATION = "C12R17.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_1a = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_1b = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1.init_1c = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .PCK_LOCATION = "C18R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26] .always_en = 1;
LUT6 ii2855 (
	. xy ( \ii2855|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[7]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2854|xy_net  )
);
defparam ii2855.PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.lut_0";
defparam ii2855.PCK_LOCATION = "C14R10.lp0.lut_0";
defparam ii2855.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
LUT6 ii2856 (
	. xy ( \ii2856|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2856.PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.lut_0";
defparam ii2856.PCK_LOCATION = "C10R9.lp0.lut_0";
defparam ii2856.config_data = 64'b1111010110110001111001001010000011110101101100011110010010100000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .PCK_LOCATION = "C16R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5] .always_en = 1;
LUT6 ii2857 (
	. xy ( \ii2857|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2857.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2857.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2857.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1]|qx_net  ),
	. di ( \ii2472|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .PCK_LOCATION = "C6R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[1] .always_en = 1;
LUT6 ii2858 (
	. xy ( \ii2858|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0]|qx_net  )
);
defparam ii2858.PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.lut_0";
defparam ii2858.PCK_LOCATION = "C14R9.lp0.lut_0";
defparam ii2858.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
REG \mcu_arbiter_func_reg[5]  (
	. qx ( \mcu_arbiter_func_reg[5]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[5] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[5] .init = 0;
defparam \mcu_arbiter_func_reg[5] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[5] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[5] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[5] .no_sr = 0;
defparam \mcu_arbiter_func_reg[5] .sr_value = 0;
defparam \mcu_arbiter_func_reg[5] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_func_reg[5] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[5] .en_inv = 0;
defparam \mcu_arbiter_func_reg[5] .always_en = 0;
LUT6 ii2860 (
	. xy ( \ii2860|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2860.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2860.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2860.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2859 (
	. xy ( \ii2859|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2858|xy_net  ),
	. f1 ( \ii2857|xy_net  ),
	. f0 ( \ii2856|xy_net  )
);
defparam ii2859.PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.lut_0";
defparam ii2859.PCK_LOCATION = "C14R9.lp0.lut_0";
defparam ii2859.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg|qx_net  ),
	. di ( \ii2075|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.PCK_LOCATION = "C14R29.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[27]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[27]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[27] .always_en = 1;
LUT6 ii2861 (
	. xy ( \ii2861|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2861.PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.lut_0";
defparam ii2861.PCK_LOCATION = "C14R9.lp0.lut_0";
defparam ii2861.config_data = 64'b1111010110110001111001001010000011110101101100011110010010100000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. di ( \ii2788|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .PCK_LOCATION = "C8R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44] .always_en = 1;
LUT6 ii2862 (
	. xy ( \ii2862|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1]|qx_net  )
);
defparam ii2862.PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.lut_0";
defparam ii2862.PCK_LOCATION = "C14R10.lp0.lut_0";
defparam ii2862.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_8__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2] .always_en = 1;
LUT6 ii2863 (
	. xy ( \ii2863|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2862|xy_net  ),
	. f1 ( \ii2861|xy_net  ),
	. f0 ( \ii2860|xy_net  )
);
defparam ii2863.PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.lut_0";
defparam ii2863.PCK_LOCATION = "C10R9.lp0.lut_0";
defparam ii2863.config_data = 64'b1111000010101010110011001100110011110000101010101100110011001100;
LUT6 ii2864 (
	. xy ( \ii2864|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2864.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2864.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2864.config_data = 64'b1111111010111010011101100011001011011100100110000101010000010000;
LUT6 ii1982_dup (
	. xy ( \ii1982_dup|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \rstn_r_reg|qx_net  ),
	. f0 ( \io_phone_rst_inst|f_id[0]_net  )
);
defparam ii1982_dup.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii1982_dup.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii1982_dup.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27] .always_en = 1;
LUT6 ii2865 (
	. xy ( \ii2865|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2864|xy_net  )
);
defparam ii2865.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2865.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2865.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2866 (
	. xy ( \ii2866|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2866.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam ii2866.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam ii2866.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2867 (
	. xy ( \ii2867|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2866|xy_net  )
);
defparam ii2867.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2867.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2867.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2]|qx_net  ),
	. di ( \ii2473|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[2] .always_en = 1;
LUT6 ii2868 (
	. xy ( \ii2868|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2868.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam ii2868.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam ii2868.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
REG \mcu_arbiter_func_reg[6]  (
	. qx ( \mcu_arbiter_func_reg[6]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[6] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[6] .init = 0;
defparam \mcu_arbiter_func_reg[6] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[6] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[6] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[6] .no_sr = 0;
defparam \mcu_arbiter_func_reg[6] .sr_value = 0;
defparam \mcu_arbiter_func_reg[6] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_func_reg[6] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[6] .en_inv = 0;
defparam \mcu_arbiter_func_reg[6] .always_en = 0;
LUT6 ii2870 (
	. xy ( \ii2870|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2870.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam ii2870.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam ii2870.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2869 (
	. xy ( \ii2869|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2868|xy_net  )
);
defparam ii2869.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2869.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2869.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[28]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[28]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[28] .always_en = 1;
LUT6 ii2871 (
	. xy ( \ii2871|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2870|xy_net  )
);
defparam ii2871.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2871.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2871.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. di ( \ii2793|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45] .always_en = 1;
LUT6 ii2872 (
	. xy ( \ii2872|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2872.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam ii2872.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam ii2872.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_8__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3] .always_en = 1;
LUT6 ii2873 (
	. xy ( \ii2873|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2872|xy_net  )
);
defparam ii2873.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2873.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2873.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2874 (
	. xy ( \ii2874|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2874.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam ii2874.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam ii2874.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[15]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2875 (
	. xy ( \ii2875|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2874|xy_net  )
);
defparam ii2875.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2875.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2875.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2876 (
	. xy ( \ii2876|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2876.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2876.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2876.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
LUT6 ii2877 (
	. xy ( \ii2877|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2876|xy_net  )
);
defparam ii2877.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2877.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2877.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3]|qx_net  ),
	. di ( \ii2474|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[3] .always_en = 1;
LUT6 ii2878 (
	. xy ( \ii2878|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2878.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2878.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2878.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
REG \mcu_arbiter_func_reg[7]  (
	. qx ( \mcu_arbiter_func_reg[7]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3321|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_func_reg[7] .latch_mode = 0;
defparam \mcu_arbiter_func_reg[7] .init = 0;
defparam \mcu_arbiter_func_reg[7] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_func_reg[7] .sr_inv = 1;
defparam \mcu_arbiter_func_reg[7] .sync_mode = 0;
defparam \mcu_arbiter_func_reg[7] .no_sr = 0;
defparam \mcu_arbiter_func_reg[7] .sr_value = 0;
defparam \mcu_arbiter_func_reg[7] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_func_reg[7] .clk_inv = 0;
defparam \mcu_arbiter_func_reg[7] .en_inv = 0;
defparam \mcu_arbiter_func_reg[7] .always_en = 0;
LUT6 ii2880 (
	. xy ( \ii2880|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2880.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii2880.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii2880.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2879 (
	. xy ( \ii2879|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2878|xy_net  )
);
defparam ii2879.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2879.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2879.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[29]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[29]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[30]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[30]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[30] .always_en = 1;
LUT6 ii2881 (
	. xy ( \ii2881|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2880|xy_net  )
);
defparam ii2881.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2881.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2881.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. di ( \ii2798|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46] .always_en = 1;
SIO io_swire_inst (
	. f_id ( )
,
	. clk_en ( ),
	. fclk ( ),
	. od ( )
,
	. oen ( ),
	. rstn ( ),
	. setn ( ),
	. PAD ( swire )
);
defparam io_swire_inst.DDR_PREG_EN = 0;
defparam io_swire_inst.FCLK_GATE_EN = 0;
defparam io_swire_inst.FOEN_SEL = 0;
defparam io_swire_inst.RSTN_SYNC = 0;
defparam io_swire_inst.OUT_SEL = 0;
defparam io_swire_inst.DDR_EN = 0;
defparam io_swire_inst.NDR = 15;
defparam io_swire_inst.VPCI_EN = 0;
defparam io_swire_inst.ID_RSTN_EN = 0;
defparam io_swire_inst.KEEP = 0;
defparam io_swire_inst.PDR = 15;
defparam io_swire_inst.SETN_INV = 0;
defparam io_swire_inst.SETN_SYNC = 0;
defparam io_swire_inst.FIN_SEL = 0;
defparam io_swire_inst.ID_SETN_EN = 0;
defparam io_swire_inst.DDR_REG_EN = 0;
defparam io_swire_inst.FOUT_SEL = 0;
defparam io_swire_inst.OEN_RSTN_EN = 0;
defparam io_swire_inst.NS_LV = 3;
defparam io_swire_inst.optional_function = "";
defparam io_swire_inst.OD_RSTN_EN = 0;
defparam io_swire_inst.RSTN_INV = 0;
defparam io_swire_inst.is_clk_io = "false";
defparam io_swire_inst.PLACE_LOCATION = "C24R5.io_guts.iob_ck.I0.I60.Iioc0";
defparam io_swire_inst.OEN_SETN_EN = 0;
defparam io_swire_inst.OEN_SEL = 1;
defparam io_swire_inst.PCK_LOCATION = "NONE";
defparam io_swire_inst.OD_SETN_EN = 0;
defparam io_swire_inst.CLK_INV = 0;
defparam io_swire_inst.is_signal_monitor_io = 1'b0;
defparam io_swire_inst.DDR_NREG_EN = 0;
defparam io_swire_inst.RX_DIG_EN = 0;
LUT6 ii2882 (
	. xy ( \ii2882|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2882.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam ii2882.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam ii2882.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_8__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4] .always_en = 1;
LUT6 ii2883 (
	. xy ( \ii2883|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2882|xy_net  )
);
defparam ii2883.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2883.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2883.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2884 (
	. xy ( \ii2884|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2884.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii2884.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii2884.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[10] .always_en = 1;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. di ( \ii2146|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.PCK_LOCATION = "C14R21.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30] .always_en = 1;
LUT6 ii2885 (
	. xy ( \ii2885|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2884|xy_net  )
);
defparam ii2885.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2885.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2885.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2886 (
	. xy ( \ii2886|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2886.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2886.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2886.config_data = 64'b1111101111101010011100110110001011011001110010000101000101000000;
LUT6 ii2887 (
	. xy ( \ii2887|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2886|xy_net  )
);
defparam ii2887.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2887.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2887.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4]|qx_net  ),
	. di ( \ii2475|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[4] .always_en = 1;
LUT6 ii2888 (
	. xy ( \ii2888|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2888.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam ii2888.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam ii2888.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2900 (
	. xy ( \ii2900|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[42]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[34]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2900.PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.lut_0";
defparam ii2900.PCK_LOCATION = "C8R16.lp0.lut_0";
defparam ii2900.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
LUT6 ii2890 (
	. xy ( \ii2890|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2890.PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.lut_0";
defparam ii2890.PCK_LOCATION = "C10R16.lp0.lut_0";
defparam ii2890.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
LUT6 ii2889 (
	. xy ( \ii2889|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2888|xy_net  )
);
defparam ii2889.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2889.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2889.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[31]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[31]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .PCK_LOCATION = "C6R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[31] .always_en = 1;
LUT6 ii2901 (
	. xy ( \ii2901|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2900|xy_net  )
);
defparam ii2901.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2901.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2901.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
LUT6 ii2891 (
	. xy ( \ii2891|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2890|xy_net  )
);
defparam ii2891.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2891.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2891.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. di ( \ii2803|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47] .always_en = 1;
REG mcu_arbiter_fifo_clr_s_reg (
	. qx ( \mcu_arbiter_fifo_clr_s_reg|qx_net  ),
	. di ( \mcu_arbiter_fifo_clr_f_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_fifo_clr_s_reg.latch_mode = 0;
defparam mcu_arbiter_fifo_clr_s_reg.init = 0;
defparam mcu_arbiter_fifo_clr_s_reg.PLACE_LOCATION = "C4R22.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_fifo_clr_s_reg.sr_inv = 1;
defparam mcu_arbiter_fifo_clr_s_reg.sync_mode = 0;
defparam mcu_arbiter_fifo_clr_s_reg.no_sr = 0;
defparam mcu_arbiter_fifo_clr_s_reg.sr_value = 0;
defparam mcu_arbiter_fifo_clr_s_reg.PCK_LOCATION = "C4R22.lp0.reg0";
defparam mcu_arbiter_fifo_clr_s_reg.clk_inv = 0;
defparam mcu_arbiter_fifo_clr_s_reg.en_inv = 0;
defparam mcu_arbiter_fifo_clr_s_reg.always_en = 1;
LUT6 ii2902 (
	. xy ( \ii2902|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[43]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[35]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2902.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii2902.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii2902.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
LUT6 ii2892 (
	. xy ( \ii2892|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2892.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2892.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2892.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_8__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5] .always_en = 1;
LUT6 ii2903 (
	. xy ( \ii2903|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2902|xy_net  )
);
defparam ii2903.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2903.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2903.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
LUT6 ii2893 (
	. xy ( \ii2893|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2892|xy_net  )
);
defparam ii2893.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2893.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2893.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
OSCV1 u_osc (
	. OSC ( \u_osc|OSC_net  )
);
defparam u_osc.osc_pd = 0;
defparam u_osc.PLACE_LOCATION = "C23R26.OSCV1";
defparam u_osc.osc_stb = 0;
defparam u_osc.PCK_LOCATION = "NONE";
LUT6 ii2904 (
	. xy ( \ii2904|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[44]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[36]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2904.PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.lut_0";
defparam ii2904.PCK_LOCATION = "C8R16.lp0.lut_0";
defparam ii2904.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2894 (
	. xy ( \ii2894|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2894.PLACE_LOCATION = "C14R15.le_tile.le_guts.lp0.lut_0";
defparam ii2894.PCK_LOCATION = "C14R15.lp0.lut_0";
defparam ii2894.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .PCK_LOCATION = "C10R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[11] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u0_hardfifo_u_inst|dout[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31] .always_en = 1;
LUT6 ii2905 (
	. xy ( \ii2905|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2904|xy_net  )
);
defparam ii2905.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.lut_0";
defparam ii2905.PCK_LOCATION = "C8R20.lp0.lut_0";
defparam ii2905.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2895 (
	. xy ( \ii2895|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2894|xy_net  )
);
defparam ii2895.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2895.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2895.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
ADD1_A carry_12_2__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_12_2__ADD_0|co_net  ),
	. s ( )
);
defparam carry_12_2__ADD_0.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_0.a_inv = "false";
defparam carry_12_2__ADD_0.PCK_LOCATION = "C16R4.lp0.add2.add0";
LUT6 ii2906 (
	. xy ( \ii2906|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[45]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[37]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2906.PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.lut_0";
defparam ii2906.PCK_LOCATION = "C8R16.lp0.lut_0";
defparam ii2906.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2896 (
	. xy ( \ii2896|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[40]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2896.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2896.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2896.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
ADD1_A carry_12_2__ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1]|qx_net  ),
	. ci ( \carry_12_2__ADD_0|co_net  ),
	. co ( \carry_12_2__ADD_1|co_net  ),
	. s ( \carry_12_2__ADD_1|s_net  )
);
defparam carry_12_2__ADD_1.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_1.a_inv = "false";
defparam carry_12_2__ADD_1.PCK_LOCATION = "C16R4.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0]|qx_net  ),
	. di ( \ii2253|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .PCK_LOCATION = "C14R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0] .always_en = 0;
LUT6 ii2907 (
	. xy ( \ii2907|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2906|xy_net  )
);
defparam ii2907.PLACE_LOCATION = "C8R21.le_tile.le_guts.lp0.lut_0";
defparam ii2907.PCK_LOCATION = "C8R21.lp0.lut_0";
defparam ii2907.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2897 (
	. xy ( \ii2897|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2896|xy_net  )
);
defparam ii2897.PLACE_LOCATION = "C10R21.le_tile.le_guts.lp0.lut_0";
defparam ii2897.PCK_LOCATION = "C10R21.lp0.lut_0";
defparam ii2897.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
ADD1_A carry_12_2__ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2]|qx_net  ),
	. ci ( \carry_12_2__ADD_1|co_net  ),
	. co ( \carry_12_2__ADD_2|co_net  ),
	. s ( \carry_12_2__ADD_2|s_net  )
);
defparam carry_12_2__ADD_2.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_2.a_inv = "false";
defparam carry_12_2__ADD_2.PCK_LOCATION = "C16R4.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5]|qx_net  ),
	. di ( \ii2476|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[5] .always_en = 1;
LUT6 ii2908 (
	. xy ( \ii2908|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2908.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam ii2908.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam ii2908.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
LUT6 ii2898 (
	. xy ( \ii2898|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[41]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2898.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam ii2898.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam ii2898.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
ADD1_A carry_12_2__ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3]|qx_net  ),
	. ci ( \carry_12_2__ADD_2|co_net  ),
	. co ( \carry_12_2__ADD_3|co_net  ),
	. s ( \carry_12_2__ADD_3|s_net  )
);
defparam carry_12_2__ADD_3.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_3.a_inv = "false";
defparam carry_12_2__ADD_3.PCK_LOCATION = "C16R4.lp0.add2.add0";
LUT6 ii2910 (
	. xy ( \ii2910|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[46]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[38]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2910.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2910.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2910.config_data = 64'b1111111011011100101110101001100001110110010101000011001000010000;
LUT6 ii2909 (
	. xy ( \ii2909|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2908|xy_net  )
);
defparam ii2909.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2909.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2909.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2899 (
	. xy ( \ii2899|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2898|xy_net  )
);
defparam ii2899.PLACE_LOCATION = "C8R21.le_tile.le_guts.lp0.lut_0";
defparam ii2899.PCK_LOCATION = "C8R21.lp0.lut_0";
defparam ii2899.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[1] .always_en = 1;
ADD1_A carry_12_2__ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4]|qx_net  ),
	. ci ( \carry_12_2__ADD_3|co_net  ),
	. co ( \carry_12_2__ADD_4|co_net  ),
	. s ( \carry_12_2__ADD_4|s_net  )
);
defparam carry_12_2__ADD_4.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_4.a_inv = "false";
defparam carry_12_2__ADD_4.PCK_LOCATION = "C16R4.lp0.add2.add0";
LUT6 ii2911 (
	. xy ( \ii2911|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2910|xy_net  )
);
defparam ii2911.PLACE_LOCATION = "C8R21.le_tile.le_guts.lp0.lut_0";
defparam ii2911.PCK_LOCATION = "C8R21.lp0.lut_0";
defparam ii2911.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48]|qx_net  ),
	. di ( \ii2808|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[48] .always_en = 1;
ADD1_A carry_12_2__ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5]|qx_net  ),
	. ci ( \carry_12_2__ADD_4|co_net  ),
	. co ( \carry_12_2__ADD_5|co_net  ),
	. s ( \carry_12_2__ADD_5|s_net  )
);
defparam carry_12_2__ADD_5.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_5.a_inv = "false";
defparam carry_12_2__ADD_5.PCK_LOCATION = "C16R4.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0]|qx_net  ),
	. di ( \ii2447|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0] .always_en = 1;
LUT6 ii2912 (
	. xy ( \ii2912|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[47]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[39]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2912.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2912.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2912.config_data = 64'b0000000100100011010001010110011110001001101010111100110111101111;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_8__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6] .always_en = 1;
ADD1_A carry_12_2__ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6]|qx_net  ),
	. ci ( \carry_12_2__ADD_5|co_net  ),
	. co ( \carry_12_2__ADD_6|co_net  ),
	. s ( \carry_12_2__ADD_6|s_net  )
);
defparam carry_12_2__ADD_6.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_6.a_inv = "false";
defparam carry_12_2__ADD_6.PCK_LOCATION = "C16R4.lp0.add2.add0";
LUT6 ii2913 (
	. xy ( \ii2913|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2912|xy_net  )
);
defparam ii2913.PLACE_LOCATION = "C10R21.le_tile.le_guts.lp0.lut_0";
defparam ii2913.PCK_LOCATION = "C10R21.lp0.lut_0";
defparam ii2913.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
ADD1_A carry_12_2__ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7]|qx_net  ),
	. ci ( \carry_12_2__ADD_6|co_net  ),
	. co ( \carry_12_2__ADD_7|co_net  ),
	. s ( \carry_12_2__ADD_7|s_net  )
);
defparam carry_12_2__ADD_7.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_7.a_inv = "false";
defparam carry_12_2__ADD_7.PCK_LOCATION = "C16R4.lp0.add2.add0";
LUT6 ii2914 (
	. xy ( \ii2914|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2914.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2914.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2914.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .PCK_LOCATION = "C10R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[12] .always_en = 1;
ADD1_A carry_12_2__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8]|qx_net  ),
	. ci ( \carry_12_2__ADD_7|co_net  ),
	. co ( \carry_12_2__ADD_8|co_net  ),
	. s ( \carry_12_2__ADD_8|s_net  )
);
defparam carry_12_2__ADD_8.PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_8.a_inv = "false";
defparam carry_12_2__ADD_8.PCK_LOCATION = "C16R5.lp0.add2.add0";
LUT6 ii2915 (
	. xy ( \ii2915|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2914|xy_net  )
);
defparam ii2915.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2915.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2915.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
ADD1_A carry_12_2__ADD_9 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9]|qx_net  ),
	. ci ( \carry_12_2__ADD_8|co_net  ),
	. co ( \carry_12_2__ADD_9|co_net  ),
	. s ( \carry_12_2__ADD_9|s_net  )
);
defparam carry_12_2__ADD_9.PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_9.a_inv = "false";
defparam carry_12_2__ADD_9.PCK_LOCATION = "C16R5.lp0.add2.add0";
LUT6 ii2916 (
	. xy ( \ii2916|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2916.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2916.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2916.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1]|qx_net  ),
	. di ( \ii2283|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0] .always_en = 1;
LUT6 ii2917 (
	. xy ( \ii2917|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2916|xy_net  )
);
defparam ii2917.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2917.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2917.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6]|qx_net  ),
	. di ( \ii2477|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[6] .always_en = 1;
LUT6 ii2918 (
	. xy ( \ii2918|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[29]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2918.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2918.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2918.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0]|qx_net  ),
	. di ( \ii2151|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0] .always_en = 0;
LUT6 ii2920 (
	. xy ( \ii2920|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[30]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2920.PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.lut_0";
defparam ii2920.PCK_LOCATION = "C10R14.lp0.lut_0";
defparam ii2920.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
LUT6 ii2919 (
	. xy ( \ii2919|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2918|xy_net  )
);
defparam ii2919.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2919.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2919.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[10] .always_en = 1;
REG \glue_dnum_s_reg[0]  (
	. qx ( \glue_dnum_s_reg[0]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[0] .latch_mode = 0;
defparam \glue_dnum_s_reg[0] .init = 0;
defparam \glue_dnum_s_reg[0] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[0] .sr_inv = 1;
defparam \glue_dnum_s_reg[0] .sync_mode = 0;
defparam \glue_dnum_s_reg[0] .no_sr = 0;
defparam \glue_dnum_s_reg[0] .sr_value = 0;
defparam \glue_dnum_s_reg[0] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[0] .clk_inv = 0;
defparam \glue_dnum_s_reg[0] .en_inv = 0;
defparam \glue_dnum_s_reg[0] .always_en = 0;
LUT6 ii3021 (
	. xy ( \ii3021|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_13__ADD_8|co_net  )
);
defparam ii3021.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.lut_0";
defparam ii3021.PCK_LOCATION = "C18R15.lp0.lut_0";
defparam ii3021.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 ii2921 (
	. xy ( \ii2921|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2920|xy_net  )
);
defparam ii2921.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2921.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2921.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50]|qx_net  ),
	. di ( \ii2821|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[50] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49]|qx_net  ),
	. di ( \ii2813|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[49] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1]|qx_net  ),
	. di ( \ii2448|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1] .always_en = 1;
LUT6 ii2922 (
	. xy ( \ii2922|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[31]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2922.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam ii2922.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam ii2922.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_8__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7] .always_en = 1;
LUT6 ii2923 (
	. xy ( \ii2923|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2922|xy_net  )
);
defparam ii2923.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2923.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2923.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
LUT6 ii2924 (
	. xy ( \ii2924|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[32]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2924.PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.lut_0";
defparam ii2924.PCK_LOCATION = "C14R14.lp0.lut_0";
defparam ii2924.config_data = 64'b0000001001000110100010101100111000010011010101111001101111011111;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[13] .always_en = 1;
LUT6 ii2925 (
	. xy ( \ii2925|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2924|xy_net  )
);
defparam ii2925.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2925.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2925.config_data = 64'b1101011100010100110101110001010011010111000101001101011100010100;
REG uut_dataReadBack_mipi_periph_dphy_direction_d_reg (
	. qx ( \uut_dataReadBack_mipi_periph_dphy_direction_d_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_dphy_direction_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.latch_mode = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.init = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.sr_inv = 1;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.sync_mode = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.no_sr = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.sr_value = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.PCK_LOCATION = "C4R8.lp0.reg0";
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.clk_inv = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.en_inv = 0;
defparam uut_dataReadBack_mipi_periph_dphy_direction_d_reg.always_en = 1;
LUT6 ii2926 (
	. xy ( \ii2926|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[33]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  )
);
defparam ii2926.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2926.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2926.config_data = 64'b1111110110111001011101010011000111101100101010000110010000100000;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc267 ,
		/* a_mac_out [23] (nc) */ nc268 ,
		/* a_mac_out [22] (nc) */ nc269 ,
		/* a_mac_out [21] (nc) */ nc270 ,
		/* a_mac_out [20] (nc) */ nc271 ,
		/* a_mac_out [19] (nc) */ nc272 ,
		/* a_mac_out [18] (nc) */ nc273 ,
		/* a_mac_out [17] (nc) */ nc274 ,
		/* a_mac_out [16] (nc) */ nc275 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc276 ,
		/* a_mac_out [2] (nc) */ nc277 ,
		/* a_mac_out [1] (nc) */ nc278 ,
		/* a_mac_out [0] (nc) */ nc279 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.PLACE_LOCATION = "C22R3.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.PCK_LOCATION = "C22R3.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2]|qx_net  ),
	. di ( \ii2284|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1] .always_en = 1;
LUT6 ii2927 (
	. xy ( \ii2927|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f0 ( \ii2926|xy_net  )
);
defparam ii2927.PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.lut_0";
defparam ii2927.PCK_LOCATION = "C10R20.lp0.lut_0";
defparam ii2927.config_data = 64'b1110101100101000111010110010100011101011001010001110101100101000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7]|qx_net  ),
	. di ( \ii2478|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_3_reg[7] .always_en = 1;
LUT6 ii2928 (
	. xy ( \ii2928|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t86_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  )
);
defparam ii2928.PLACE_LOCATION = "C6R21.le_tile.le_guts.lp0.lut_0";
defparam ii2928.PCK_LOCATION = "C6R21.lp0.lut_0";
defparam ii2928.config_data = 64'b0110000001100000011000000110000001100000011000000110000001100000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1]|qx_net  ),
	. di ( \ii2165|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1] .always_en = 0;
LUT6 ii2930 (
	. xy ( \ii2930|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[25]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[1]_net  )
);
defparam ii2930.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2930.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2930.config_data = 64'b1010111111001111101000001100000010101111110011111010000011000000;
LUT6 ii2929 (
	. xy ( \ii2929|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[24]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[0]_net  )
);
defparam ii2929.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2929.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2929.config_data = 64'b1010111111001111101000001100000010101111110011111010000011000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .PCK_LOCATION = "C18R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .PCK_LOCATION = "C8R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[11] .always_en = 1;
REG \glue_dnum_s_reg[1]  (
	. qx ( \glue_dnum_s_reg[1]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[1] .latch_mode = 0;
defparam \glue_dnum_s_reg[1] .init = 0;
defparam \glue_dnum_s_reg[1] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[1] .sr_inv = 1;
defparam \glue_dnum_s_reg[1] .sync_mode = 0;
defparam \glue_dnum_s_reg[1] .no_sr = 0;
defparam \glue_dnum_s_reg[1] .sr_value = 0;
defparam \glue_dnum_s_reg[1] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[1] .clk_inv = 0;
defparam \glue_dnum_s_reg[1] .en_inv = 0;
defparam \glue_dnum_s_reg[1] .always_en = 0;
LUT6 ii2931 (
	. xy ( \ii2931|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[2]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[26]_net  )
);
defparam ii2931.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2931.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2931.config_data = 64'b1100111110101111110000001010000011001111101011111100000010100000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51]|qx_net  ),
	. di ( \ii2826|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[51] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2]|qx_net  ),
	. di ( \ii2449|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .PCK_LOCATION = "C10R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0] .always_en = 1;
LUT6 ii2932 (
	. xy ( \ii2932|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[3]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[27]_net  )
);
defparam ii2932.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2932.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2932.config_data = 64'b1100111110101111110000001010000011001111101011111100000010100000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net  ),
	. di ( \ii3195|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .PCK_LOCATION = "C20R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8] .always_en = 1;
FIFO18K glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst (
	. dout ( {
		/* dout [63] (nc) */ nc280 ,
		/* dout [62] (nc) */ nc281 ,
		/* dout [61] (nc) */ nc282 ,
		/* dout [60] (nc) */ nc283 ,
		/* dout [59] (nc) */ nc284 ,
		/* dout [58] (nc) */ nc285 ,
		/* dout [57] (nc) */ nc286 ,
		/* dout [56] (nc) */ nc287 ,
		/* dout [55] (nc) */ nc288 ,
		/* dout [54] (nc) */ nc289 ,
		/* dout [53] (nc) */ nc290 ,
		/* dout [52] (nc) */ nc291 ,
		/* dout [51] (nc) */ nc292 ,
		/* dout [50] (nc) */ nc293 ,
		/* dout [49] (nc) */ nc294 ,
		/* dout [48] (nc) */ nc295 ,
		/* dout [47] (nc) */ nc296 ,
		/* dout [46] (nc) */ nc297 ,
		/* dout [45] (nc) */ nc298 ,
		/* dout [44] (nc) */ nc299 ,
		/* dout [43] (nc) */ nc300 ,
		/* dout [42] (nc) */ nc301 ,
		/* dout [41] (nc) */ nc302 ,
		/* dout [40] (nc) */ nc303 ,
		/* dout [39] (nc) */ nc304 ,
		/* dout [38] (nc) */ nc305 ,
		/* dout [37] (nc) */ nc306 ,
		/* dout [36] (nc) */ nc307 ,
		/* dout [35] (nc) */ nc308 ,
		/* dout [34] (nc) */ nc309 ,
		/* dout [33] (nc) */ nc310 ,
		/* dout [32] (nc) */ nc311 ,
		/* dout [31] (nc) */ nc312 ,
		/* dout [30] (nc) */ nc313 ,
		/* dout [29] (nc) */ nc314 ,
		/* dout [28] (nc) */ nc315 ,
		/* dout [27] (nc) */ nc316 ,
		/* dout [26] (nc) */ nc317 ,
		/* dout [25] (nc) */ nc318 ,
		/* dout [24] (nc) */ nc319 ,
		/* dout [23] (nc) */ nc320 ,
		/* dout [22] (nc) */ nc321 ,
		/* dout [21] (nc) */ nc322 ,
		/* dout [20] (nc) */ nc323 ,
		/* dout [19] (nc) */ nc324 ,
		/* dout [18] (nc) */ nc325 ,
		/* dout [17] (nc) */ nc326 ,
		/* dout [16] (nc) */ nc327 ,
		/* dout [15] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[15]_net ,
		/* dout [14] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[14]_net ,
		/* dout [13] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[13]_net ,
		/* dout [12] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[12]_net ,
		/* dout [11] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[11]_net ,
		/* dout [10] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[10]_net ,
		/* dout [9] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[9]_net ,
		/* dout [8] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[8]_net ,
		/* dout [7] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[7]_net ,
		/* dout [6] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[6]_net ,
		/* dout [5] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[5]_net ,
		/* dout [4] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[4]_net ,
		/* dout [3] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[3]_net ,
		/* dout [2] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[2]_net ,
		/* dout [1] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[1]_net ,
		/* dout [0] */ \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[0]_net 
	} ),
	. doutp ( )
,
	. din ( {
		/* din [63] */ \GND_0_inst|Y_net ,
		/* din [62] */ \GND_0_inst|Y_net ,
		/* din [61] */ \GND_0_inst|Y_net ,
		/* din [60] */ \GND_0_inst|Y_net ,
		/* din [59] */ \GND_0_inst|Y_net ,
		/* din [58] */ \GND_0_inst|Y_net ,
		/* din [57] */ \GND_0_inst|Y_net ,
		/* din [56] */ \GND_0_inst|Y_net ,
		/* din [55] */ \GND_0_inst|Y_net ,
		/* din [54] */ \GND_0_inst|Y_net ,
		/* din [53] */ \GND_0_inst|Y_net ,
		/* din [52] */ \GND_0_inst|Y_net ,
		/* din [51] */ \GND_0_inst|Y_net ,
		/* din [50] */ \GND_0_inst|Y_net ,
		/* din [49] */ \GND_0_inst|Y_net ,
		/* din [48] */ \GND_0_inst|Y_net ,
		/* din [47] */ \GND_0_inst|Y_net ,
		/* din [46] */ \GND_0_inst|Y_net ,
		/* din [45] */ \GND_0_inst|Y_net ,
		/* din [44] */ \GND_0_inst|Y_net ,
		/* din [43] */ \GND_0_inst|Y_net ,
		/* din [42] */ \GND_0_inst|Y_net ,
		/* din [41] */ \GND_0_inst|Y_net ,
		/* din [40] */ \GND_0_inst|Y_net ,
		/* din [39] */ \GND_0_inst|Y_net ,
		/* din [38] */ \GND_0_inst|Y_net ,
		/* din [37] */ \GND_0_inst|Y_net ,
		/* din [36] */ \GND_0_inst|Y_net ,
		/* din [35] */ \GND_0_inst|Y_net ,
		/* din [34] */ \GND_0_inst|Y_net ,
		/* din [33] */ \GND_0_inst|Y_net ,
		/* din [32] */ \GND_0_inst|Y_net ,
		/* din [31] */ \GND_0_inst|Y_net ,
		/* din [30] */ \GND_0_inst|Y_net ,
		/* din [29] */ \GND_0_inst|Y_net ,
		/* din [28] */ \GND_0_inst|Y_net ,
		/* din [27] */ \GND_0_inst|Y_net ,
		/* din [26] */ \GND_0_inst|Y_net ,
		/* din [25] */ \GND_0_inst|Y_net ,
		/* din [24] */ \GND_0_inst|Y_net ,
		/* din [23] */ \GND_0_inst|Y_net ,
		/* din [22] */ \GND_0_inst|Y_net ,
		/* din [21] */ \GND_0_inst|Y_net ,
		/* din [20] */ \GND_0_inst|Y_net ,
		/* din [19] */ \GND_0_inst|Y_net ,
		/* din [18] */ \GND_0_inst|Y_net ,
		/* din [17] */ \GND_0_inst|Y_net ,
		/* din [16] */ \GND_0_inst|Y_net ,
		/* din [15] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7]|qx_net ,
		/* din [14] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6]|qx_net ,
		/* din [13] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5]|qx_net ,
		/* din [12] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4]|qx_net ,
		/* din [11] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3]|qx_net ,
		/* din [10] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2]|qx_net ,
		/* din [9] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1]|qx_net ,
		/* din [8] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0]|qx_net ,
		/* din [7] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15]|qx_net ,
		/* din [6] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14]|qx_net ,
		/* din [5] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13]|qx_net ,
		/* din [4] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12]|qx_net ,
		/* din [3] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11]|qx_net ,
		/* din [2] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10]|qx_net ,
		/* din [1] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9]|qx_net ,
		/* din [0] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8]|qx_net 
	} ),
	. dinp ( {
		/* dinp [7] */ \GND_0_inst|Y_net ,
		/* dinp [6] */ \GND_0_inst|Y_net ,
		/* dinp [5] */ \GND_0_inst|Y_net ,
		/* dinp [4] */ \GND_0_inst|Y_net ,
		/* dinp [3] */ \GND_0_inst|Y_net ,
		/* dinp [2] */ \GND_0_inst|Y_net ,
		/* dinp [1] */ \GND_0_inst|Y_net ,
		/* dinp [0] */ \GND_0_inst|Y_net 
	} ),
	. writeclk ( \u_pll_pll_u0|CO0_net  ),
	. readclk ( \u_gbuf_u_gbuf|out_net  ),
	. writeen ( \ii1988|xy_net  ),
	. readen ( \ii1985|xy_net  ),
	. reset ( \ii1987|xy_net  ),
	. regce ( \VCC_0_inst|Y_net  ),
	. writesave ( \GND_0_inst|Y_net  ),
	. writedrop ( \GND_0_inst|Y_net  ),
	. full ( ),
	. empty ( ),
	. almostfull ( ),
	. almostempty ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|almostempty_net  ),
	. overflow ( ),
	. underflow ( ),
	. eccoutdberr ( ),
	. eccoutsberr ( ),
	. eccreadaddr ( )
,
	. eccindberr ( \GND_0_inst|Y_net  ),
	. eccinsberr ( \GND_0_inst|Y_net  ),
	. writedropflag ( )
);
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.eccwriteen = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.writeclk_inv = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.eccreaden = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.readclk_inv = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.use_parity = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.outreg = 1;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.almostfullth = 988;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.almostemptyth = 512;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.writewidth = 18;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.readwidth = 18;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.peek = 1;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.PLACE_LOCATION = "C12R25.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst.PCK_LOCATION = "C12R25.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
LUT6 ii2933 (
	. xy ( \ii2933|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[4]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[28]_net  )
);
defparam ii2933.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2933.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2933.config_data = 64'b1100111110101111110000001010000011001111101011111100000010100000;
LUT6 ii2934 (
	. xy ( \ii2934|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[5]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[29]_net  )
);
defparam ii2934.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2934.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2934.config_data = 64'b1100111110101111110000001010000011001111101011111100000010100000;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[14] .always_en = 1;
LUT6 u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly (
	. xy ( \u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mipi_inst_u_mipi2|clk_net  )
);
defparam u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp1.lut_1";
defparam u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly.PCK_LOCATION = "NONE";
defparam u0_mipi1_clkdly_genblk1_3__u_mipi_clkdly.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3]|qx_net  ),
	. di ( \ii2285|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2]|qx_net  ),
	. di ( \ii2178|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .PCK_LOCATION = "C8R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[12] .always_en = 1;
REG \glue_dnum_s_reg[2]  (
	. qx ( \glue_dnum_s_reg[2]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[2] .latch_mode = 0;
defparam \glue_dnum_s_reg[2] .init = 0;
defparam \glue_dnum_s_reg[2] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[2] .sr_inv = 1;
defparam \glue_dnum_s_reg[2] .sync_mode = 0;
defparam \glue_dnum_s_reg[2] .no_sr = 0;
defparam \glue_dnum_s_reg[2] .sr_value = 0;
defparam \glue_dnum_s_reg[2] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[2] .clk_inv = 0;
defparam \glue_dnum_s_reg[2] .en_inv = 0;
defparam \glue_dnum_s_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52]|qx_net  ),
	. di ( \ii2831|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[52] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3]|qx_net  ),
	. di ( \ii2450|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .PCK_LOCATION = "C10R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_d_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[0]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[15] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4]|qx_net  ),
	. di ( \ii2286|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3]|qx_net  ),
	. di ( \ii2189|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1] .always_en = 1;
LUT6 ii3050 (
	. xy ( \ii3050|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_3__ADD_8|co_net  )
);
defparam ii3050.PLACE_LOCATION = "C14R6.le_tile.le_guts.lp0.lut_0";
defparam ii3050.PCK_LOCATION = "C14R6.lp0.lut_0";
defparam ii3050.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In1p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[13] .always_en = 1;
ADD1_A carry_9_13__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_13__ADD_0|co_net  ),
	. s ( \carry_9_13__ADD_0|s_net  )
);
defparam carry_9_13__ADD_0.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_0.a_inv = "true";
defparam carry_9_13__ADD_0.PCK_LOCATION = "C10R15.lp0.add2.add0";
REG \glue_dnum_s_reg[3]  (
	. qx ( \glue_dnum_s_reg[3]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[3] .latch_mode = 0;
defparam \glue_dnum_s_reg[3] .init = 0;
defparam \glue_dnum_s_reg[3] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[3] .sr_inv = 1;
defparam \glue_dnum_s_reg[3] .sync_mode = 0;
defparam \glue_dnum_s_reg[3] .no_sr = 0;
defparam \glue_dnum_s_reg[3] .sr_value = 0;
defparam \glue_dnum_s_reg[3] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[3] .clk_inv = 0;
defparam \glue_dnum_s_reg[3] .en_inv = 0;
defparam \glue_dnum_s_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53]|qx_net  ),
	. di ( \ii2836|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .PCK_LOCATION = "C10R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[53] .always_en = 1;
ADD1_A carry_9_13__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1]|qx_net  ),
	. ci ( \carry_9_13__ADD_0|co_net  ),
	. co ( \carry_9_13__ADD_1|co_net  ),
	. s ( \carry_9_13__ADD_1|s_net  )
);
defparam carry_9_13__ADD_1.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_1.a_inv = "true";
defparam carry_9_13__ADD_1.PCK_LOCATION = "C10R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4]|qx_net  ),
	. di ( \ii2451|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t71_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t71_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.PCK_LOCATION = "C20R22.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t71_out1_reg.always_en = 1;
ADD1_A carry_9_13__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2]|qx_net  ),
	. ci ( \carry_9_13__ADD_1|co_net  ),
	. co ( \carry_9_13__ADD_2|co_net  ),
	. s ( \carry_9_13__ADD_2|s_net  )
);
defparam carry_9_13__ADD_2.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_2.a_inv = "true";
defparam carry_9_13__ADD_2.PCK_LOCATION = "C10R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_rx_cmd_d_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[1]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[1] .always_en = 1;
ADD1_A carry_9_13__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3]|qx_net  ),
	. ci ( \carry_9_13__ADD_2|co_net  ),
	. co ( \carry_9_13__ADD_3|co_net  ),
	. s ( \carry_9_13__ADD_3|s_net  )
);
defparam carry_9_13__ADD_3.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_3.a_inv = "true";
defparam carry_9_13__ADD_3.PCK_LOCATION = "C10R15.lp0.add2.add0";
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc328 ,
		/* a_mac_out [23] (nc) */ nc329 ,
		/* a_mac_out [22] (nc) */ nc330 ,
		/* a_mac_out [21] (nc) */ nc331 ,
		/* a_mac_out [20] (nc) */ nc332 ,
		/* a_mac_out [19] (nc) */ nc333 ,
		/* a_mac_out [18] (nc) */ nc334 ,
		/* a_mac_out [17] (nc) */ nc335 ,
		/* a_mac_out [16] (nc) */ nc336 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc337 ,
		/* a_mac_out [2] (nc) */ nc338 ,
		/* a_mac_out [1] (nc) */ nc339 ,
		/* a_mac_out [0] (nc) */ nc340 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.PLACE_LOCATION = "C22R5.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.PCK_LOCATION = "C22R5.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[16] .always_en = 1;
ADD1_A carry_9_13__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4]|qx_net  ),
	. ci ( \carry_9_13__ADD_3|co_net  ),
	. co ( \carry_9_13__ADD_4|co_net  ),
	. s ( \carry_9_13__ADD_4|s_net  )
);
defparam carry_9_13__ADD_4.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_4.a_inv = "true";
defparam carry_9_13__ADD_4.PCK_LOCATION = "C10R15.lp0.add2.add0";
ADD1_A carry_9_13__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5]|qx_net  ),
	. ci ( \carry_9_13__ADD_4|co_net  ),
	. co ( \carry_9_13__ADD_5|co_net  ),
	. s ( \carry_9_13__ADD_5|s_net  )
);
defparam carry_9_13__ADD_5.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_5.a_inv = "true";
defparam carry_9_13__ADD_5.PCK_LOCATION = "C10R15.lp0.add2.add0";
ADD1_A carry_9_13__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6]|qx_net  ),
	. ci ( \carry_9_13__ADD_5|co_net  ),
	. co ( \carry_9_13__ADD_6|co_net  ),
	. s ( \carry_9_13__ADD_6|s_net  )
);
defparam carry_9_13__ADD_6.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_6.a_inv = "true";
defparam carry_9_13__ADD_6.PCK_LOCATION = "C10R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5]|qx_net  ),
	. di ( \ii2287|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4] .always_en = 1;
ADD1_A carry_9_13__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7]|qx_net  ),
	. ci ( \carry_9_13__ADD_6|co_net  ),
	. co ( \carry_9_13__ADD_7|co_net  ),
	. s ( \carry_9_13__ADD_7|s_net  )
);
defparam carry_9_13__ADD_7.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_7.a_inv = "true";
defparam carry_9_13__ADD_7.PCK_LOCATION = "C10R15.lp0.add2.add0";
ADD1_A carry_9_13__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_13__ADD_7|co_net  ),
	. co ( \carry_9_13__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_13__ADD_8.PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_13__ADD_8.a_inv = "false";
defparam carry_9_13__ADD_8.PCK_LOCATION = "C10R16.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4]|qx_net  ),
	. di ( \ii2200|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[14] .always_en = 1;
REG \glue_dnum_s_reg[4]  (
	. qx ( \glue_dnum_s_reg[4]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[4] .latch_mode = 0;
defparam \glue_dnum_s_reg[4] .init = 0;
defparam \glue_dnum_s_reg[4] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[4] .sr_inv = 1;
defparam \glue_dnum_s_reg[4] .sync_mode = 0;
defparam \glue_dnum_s_reg[4] .no_sr = 0;
defparam \glue_dnum_s_reg[4] .sr_value = 0;
defparam \glue_dnum_s_reg[4] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[4] .clk_inv = 0;
defparam \glue_dnum_s_reg[4] .en_inv = 0;
defparam \glue_dnum_s_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54]|qx_net  ),
	. di ( \ii2841|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[54] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5]|qx_net  ),
	. di ( \ii2452|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_d_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[2]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[2] .always_en = 1;
LUT6 ii2963 (
	. xy ( \ii2963|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_ADD_8|co_net  )
);
defparam ii2963.PLACE_LOCATION = "C14R5.le_tile.le_guts.lp0.lut_0";
defparam ii2963.PCK_LOCATION = "C14R5.lp0.lut_0";
defparam ii2963.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[17] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[7]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
ADD1_A carry_9_3__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_3__ADD_0|co_net  ),
	. s ( \carry_9_3__ADD_0|s_net  )
);
defparam carry_9_3__ADD_0.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_0.a_inv = "true";
defparam carry_9_3__ADD_0.PCK_LOCATION = "C10R12.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6]|qx_net  ),
	. di ( \ii2288|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5] .always_en = 1;
ADD1_A carry_9_3__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1]|qx_net  ),
	. ci ( \carry_9_3__ADD_0|co_net  ),
	. co ( \carry_9_3__ADD_1|co_net  ),
	. s ( \carry_9_3__ADD_1|s_net  )
);
defparam carry_9_3__ADD_1.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_1.a_inv = "true";
defparam carry_9_3__ADD_1.PCK_LOCATION = "C10R12.lp0.add2.add0";
ADD1_A carry_9_3__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2]|qx_net  ),
	. ci ( \carry_9_3__ADD_1|co_net  ),
	. co ( \carry_9_3__ADD_2|co_net  ),
	. s ( \carry_9_3__ADD_2|s_net  )
);
defparam carry_9_3__ADD_2.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_2.a_inv = "true";
defparam carry_9_3__ADD_2.PCK_LOCATION = "C10R12.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5]|qx_net  ),
	. di ( \ii2211|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[15] .always_en = 1;
ADD1_A carry_9_3__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3]|qx_net  ),
	. ci ( \carry_9_3__ADD_2|co_net  ),
	. co ( \carry_9_3__ADD_3|co_net  ),
	. s ( \carry_9_3__ADD_3|s_net  )
);
defparam carry_9_3__ADD_3.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_3.a_inv = "true";
defparam carry_9_3__ADD_3.PCK_LOCATION = "C10R12.lp0.add2.add0";
REG \glue_dnum_s_reg[5]  (
	. qx ( \glue_dnum_s_reg[5]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[5] .latch_mode = 0;
defparam \glue_dnum_s_reg[5] .init = 0;
defparam \glue_dnum_s_reg[5] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[5] .sr_inv = 1;
defparam \glue_dnum_s_reg[5] .sync_mode = 0;
defparam \glue_dnum_s_reg[5] .no_sr = 0;
defparam \glue_dnum_s_reg[5] .sr_value = 0;
defparam \glue_dnum_s_reg[5] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[5] .clk_inv = 0;
defparam \glue_dnum_s_reg[5] .en_inv = 0;
defparam \glue_dnum_s_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55]|qx_net  ),
	. di ( \ii2846|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[55] .always_en = 1;
ADD1_A carry_9_3__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4]|qx_net  ),
	. ci ( \carry_9_3__ADD_3|co_net  ),
	. co ( \carry_9_3__ADD_4|co_net  ),
	. s ( \carry_9_3__ADD_4|s_net  )
);
defparam carry_9_3__ADD_4.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_4.a_inv = "true";
defparam carry_9_3__ADD_4.PCK_LOCATION = "C10R12.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6]|qx_net  ),
	. di ( \ii2453|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[31]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf.PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf.PCK_LOCATION = "C4R11.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[2] .always_en = 1;
ADD1_A carry_9_3__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5]|qx_net  ),
	. ci ( \carry_9_3__ADD_4|co_net  ),
	. co ( \carry_9_3__ADD_5|co_net  ),
	. s ( \carry_9_3__ADD_5|s_net  )
);
defparam carry_9_3__ADD_5.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_5.a_inv = "true";
defparam carry_9_3__ADD_5.PCK_LOCATION = "C10R12.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_rx_cmd_d_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[3]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[3] .always_en = 1;
ADD1_A carry_9_3__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6]|qx_net  ),
	. ci ( \carry_9_3__ADD_5|co_net  ),
	. co ( \carry_9_3__ADD_6|co_net  ),
	. s ( \carry_9_3__ADD_6|s_net  )
);
defparam carry_9_3__ADD_6.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_6.a_inv = "true";
defparam carry_9_3__ADD_6.PCK_LOCATION = "C10R12.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[18] .always_en = 1;
ADD1_A carry_9_3__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7]|qx_net  ),
	. ci ( \carry_9_3__ADD_6|co_net  ),
	. co ( \carry_9_3__ADD_7|co_net  ),
	. s ( \carry_9_3__ADD_7|s_net  )
);
defparam carry_9_3__ADD_7.PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_7.a_inv = "true";
defparam carry_9_3__ADD_7.PCK_LOCATION = "C10R12.lp0.add2.add0";
ADD1_A carry_9_3__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_3__ADD_7|co_net  ),
	. co ( \carry_9_3__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_3__ADD_8.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_3__ADD_8.a_inv = "false";
defparam carry_9_3__ADD_8.PCK_LOCATION = "C10R13.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7]|qx_net  ),
	. di ( \ii2289|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .PLACE_LOCATION = "C6R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .PCK_LOCATION = "C6R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6]|qx_net  ),
	. di ( \ii2216|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4] .always_en = 1;
LUT6 ii3079 (
	. xy ( \ii3079|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_4__ADD_8|co_net  )
);
defparam ii3079.PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.lut_0";
defparam ii3079.PCK_LOCATION = "C10R7.lp0.lut_0";
defparam ii3079.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .PCK_LOCATION = "C4R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[16] .always_en = 1;
REG \glue_dnum_s_reg[6]  (
	. qx ( \glue_dnum_s_reg[6]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[6] .latch_mode = 0;
defparam \glue_dnum_s_reg[6] .init = 0;
defparam \glue_dnum_s_reg[6] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[6] .sr_inv = 1;
defparam \glue_dnum_s_reg[6] .sync_mode = 0;
defparam \glue_dnum_s_reg[6] .no_sr = 0;
defparam \glue_dnum_s_reg[6] .sr_value = 0;
defparam \glue_dnum_s_reg[6] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_dnum_s_reg[6] .clk_inv = 0;
defparam \glue_dnum_s_reg[6] .en_inv = 0;
defparam \glue_dnum_s_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7]|qx_net  ),
	. di ( \ii2454|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .PCK_LOCATION = "C14R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5] .always_en = 1;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc341 ,
		/* a_mac_out [23] (nc) */ nc342 ,
		/* a_mac_out [22] (nc) */ nc343 ,
		/* a_mac_out [21] (nc) */ nc344 ,
		/* a_mac_out [20] (nc) */ nc345 ,
		/* a_mac_out [19] (nc) */ nc346 ,
		/* a_mac_out [18] (nc) */ nc347 ,
		/* a_mac_out [17] (nc) */ nc348 ,
		/* a_mac_out [16] (nc) */ nc349 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc350 ,
		/* a_mac_out [2] (nc) */ nc351 ,
		/* a_mac_out [1] (nc) */ nc352 ,
		/* a_mac_out [0] (nc) */ nc353 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.PLACE_LOCATION = "C22R7.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.PCK_LOCATION = "C22R7.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_d_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[4]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[20] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8]|qx_net  ),
	. di ( \ii2290|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .PLACE_LOCATION = "C6R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .PCK_LOCATION = "C6R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7]|qx_net  ),
	. di ( \ii2217|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_4__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .PCK_LOCATION = "C4R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[17] .always_en = 1;
REG \glue_dnum_s_reg[7]  (
	. qx ( \glue_dnum_s_reg[7]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[7] .latch_mode = 0;
defparam \glue_dnum_s_reg[7] .init = 0;
defparam \glue_dnum_s_reg[7] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[7] .sr_inv = 1;
defparam \glue_dnum_s_reg[7] .sync_mode = 0;
defparam \glue_dnum_s_reg[7] .no_sr = 0;
defparam \glue_dnum_s_reg[7] .sr_value = 0;
defparam \glue_dnum_s_reg[7] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_dnum_s_reg[7] .clk_inv = 0;
defparam \glue_dnum_s_reg[7] .en_inv = 0;
defparam \glue_dnum_s_reg[7] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6] .always_en = 1;
LUT6 ii2992 (
	. xy ( \ii2992|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_12__ADD_8|co_net  )
);
defparam ii2992.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.lut_0";
defparam ii2992.PCK_LOCATION = "C18R13.lp0.lut_0";
defparam ii2992.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_d_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[5]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_d_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[21] .always_en = 1;
ADD1_A carry_12_ADD_10 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10]|qx_net  ),
	. ci ( \carry_12_ADD_9|co_net  ),
	. co ( \carry_12_ADD_10|co_net  ),
	. s ( \carry_12_ADD_10|s_net  )
);
defparam carry_12_ADD_10.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_10.a_inv = "false";
defparam carry_12_ADD_10.PCK_LOCATION = "C14R23.lp0.add2.add0";
ADD1_A carry_12_ADD_11 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11]|qx_net  ),
	. ci ( \carry_12_ADD_10|co_net  ),
	. co ( ),
	. s ( \carry_12_ADD_11|s_net  )
);
defparam carry_12_ADD_11.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_11.a_inv = "false";
defparam carry_12_ADD_11.PCK_LOCATION = "C14R23.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9]|qx_net  ),
	. di ( \ii2291|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .PLACE_LOCATION = "C8R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .PCK_LOCATION = "C8R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .PCK_LOCATION = "C4R6.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[21]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG glue_rx_packet_tx_packet_u_scaler_t36_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t36_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_out1_1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.PCK_LOCATION = "C16R14.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t36_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0] .always_en = 1;
LUT6 ii3108 (
	. xy ( \ii3108|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_5__ADD_8|co_net  )
);
defparam ii3108.PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.lut_0";
defparam ii3108.PCK_LOCATION = "C10R7.lp0.lut_0";
defparam ii3108.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8]|qx_net  ),
	. di ( \ii2218|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_4__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .PLACE_LOCATION = "C4R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .PCK_LOCATION = "C4R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[18] .always_en = 1;
REG \glue_dnum_s_reg[8]  (
	. qx ( \glue_dnum_s_reg[8]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[16]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[8] .latch_mode = 0;
defparam \glue_dnum_s_reg[8] .init = 0;
defparam \glue_dnum_s_reg[8] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[8] .sr_inv = 1;
defparam \glue_dnum_s_reg[8] .sync_mode = 0;
defparam \glue_dnum_s_reg[8] .no_sr = 0;
defparam \glue_dnum_s_reg[8] .sr_value = 0;
defparam \glue_dnum_s_reg[8] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_dnum_s_reg[8] .clk_inv = 0;
defparam \glue_dnum_s_reg[8] .en_inv = 0;
defparam \glue_dnum_s_reg[8] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In1p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[22] .always_en = 1;
REG glue_pasm_cmd_rq_o_reg (
	. qx ( \glue_pasm_cmd_rq_o_reg|qx_net  ),
	. di ( \ii2134|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_pasm_cmd_rq_o_reg.latch_mode = 0;
defparam glue_pasm_cmd_rq_o_reg.init = 0;
defparam glue_pasm_cmd_rq_o_reg.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.reg0";
defparam glue_pasm_cmd_rq_o_reg.sr_inv = 1;
defparam glue_pasm_cmd_rq_o_reg.sync_mode = 0;
defparam glue_pasm_cmd_rq_o_reg.no_sr = 0;
defparam glue_pasm_cmd_rq_o_reg.sr_value = 0;
defparam glue_pasm_cmd_rq_o_reg.PCK_LOCATION = "C14R30.lp0.reg0";
defparam glue_pasm_cmd_rq_o_reg.clk_inv = 0;
defparam glue_pasm_cmd_rq_o_reg.en_inv = 0;
defparam glue_pasm_cmd_rq_o_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .PCK_LOCATION = "C4R6.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0]|qx_net  ),
	. di ( \ii2463|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9]|qx_net  ),
	. di ( \ii2219|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7] .always_en = 1;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc354 ,
		/* a_mac_out [23] (nc) */ nc355 ,
		/* a_mac_out [22] (nc) */ nc356 ,
		/* a_mac_out [21] (nc) */ nc357 ,
		/* a_mac_out [20] (nc) */ nc358 ,
		/* a_mac_out [19] (nc) */ nc359 ,
		/* a_mac_out [18] (nc) */ nc360 ,
		/* a_mac_out [17] (nc) */ nc361 ,
		/* a_mac_out [16] (nc) */ nc362 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc363 ,
		/* a_mac_out [2] (nc) */ nc364 ,
		/* a_mac_out [1] (nc) */ nc365 ,
		/* a_mac_out [0] (nc) */ nc366 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.PLACE_LOCATION = "C22R9.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.PCK_LOCATION = "C22R9.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_4__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[20] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[19] .always_en = 1;
REG \glue_dnum_s_reg[9]  (
	. qx ( \glue_dnum_s_reg[9]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[17]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[9] .latch_mode = 0;
defparam \glue_dnum_s_reg[9] .init = 0;
defparam \glue_dnum_s_reg[9] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[9] .sr_inv = 1;
defparam \glue_dnum_s_reg[9] .sync_mode = 0;
defparam \glue_dnum_s_reg[9] .no_sr = 0;
defparam \glue_dnum_s_reg[9] .sr_value = 0;
defparam \glue_dnum_s_reg[9] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_dnum_s_reg[9] .clk_inv = 0;
defparam \glue_dnum_s_reg[9] .en_inv = 0;
defparam \glue_dnum_s_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .PLACE_LOCATION = "C8R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .PCK_LOCATION = "C8R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[23] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1]|qx_net  ),
	. di ( \ii2464|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_4__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[21] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[11]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[24] .always_en = 1;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. di ( \ii2148|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.PCK_LOCATION = "C14R22.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg.always_en = 1;
LUT6 ii3137 (
	. xy ( \ii3137|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_6__ADD_8|co_net  )
);
defparam ii3137.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii3137.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii3137.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2]|qx_net  ),
	. di ( \ii2465|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_4__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[22] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10]|qx_net  ),
	. di ( \ii2281|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[25] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0]|qx_net  ),
	. di ( \ii3374|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0] .always_en = 0;
REG glue_rx_packet_tx_packet_fifo_vs_reg (
	. qx ( \glue_rx_packet_tx_packet_fifo_vs_reg|qx_net  ),
	. di ( \ii2142|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_fifo_vs_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.init = 0;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_fifo_vs_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.sr_value = 1;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.PCK_LOCATION = "C18R14.lp0.reg0";
defparam glue_rx_packet_tx_packet_fifo_vs_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_vs_reg.always_en = 1;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc367 ,
		/* a_mac_out [23] (nc) */ nc368 ,
		/* a_mac_out [22] (nc) */ nc369 ,
		/* a_mac_out [21] (nc) */ nc370 ,
		/* a_mac_out [20] (nc) */ nc371 ,
		/* a_mac_out [19] (nc) */ nc372 ,
		/* a_mac_out [18] (nc) */ nc373 ,
		/* a_mac_out [17] (nc) */ nc374 ,
		/* a_mac_out [16] (nc) */ nc375 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc376 ,
		/* a_mac_out [2] (nc) */ nc377 ,
		/* a_mac_out [1] (nc) */ nc378 ,
		/* a_mac_out [0] (nc) */ nc379 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.PLACE_LOCATION = "C22R23.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.PCK_LOCATION = "C22R23.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3]|qx_net  ),
	. di ( \ii2466|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_4__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[23] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11]|qx_net  ),
	. di ( \ii2282|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2254|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[26] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1]|qx_net  ),
	. di ( \ii3383|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4]|qx_net  ),
	. di ( \ii2467|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_4__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[24] .always_en = 1;
REG glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg.always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[27] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2]|qx_net  ),
	. di ( \ii3371|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2] .always_en = 0;
ADD1_A carry_12_1__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_12_1__ADD_0|co_net  ),
	. s ( )
);
defparam carry_12_1__ADD_0.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_0.a_inv = "false";
defparam carry_12_1__ADD_0.PCK_LOCATION = "C18R4.lp0.add2.add0";
LUT6 ii3166 (
	. xy ( \ii3166|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_7__ADD_8|co_net  )
);
defparam ii3166.PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.lut_0";
defparam ii3166.PCK_LOCATION = "C20R17.lp0.lut_0";
defparam ii3166.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
ADD1_A carry_12_1__ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1]|qx_net  ),
	. ci ( \carry_12_1__ADD_0|co_net  ),
	. co ( \carry_12_1__ADD_1|co_net  ),
	. s ( \carry_12_1__ADD_1|s_net  )
);
defparam carry_12_1__ADD_1.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_1.a_inv = "false";
defparam carry_12_1__ADD_1.PCK_LOCATION = "C18R4.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[4] .always_en = 1;
ADD1_A carry_12_1__ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2]|qx_net  ),
	. ci ( \carry_12_1__ADD_1|co_net  ),
	. co ( \carry_12_1__ADD_2|co_net  ),
	. s ( \carry_12_1__ADD_2|s_net  )
);
defparam carry_12_1__ADD_2.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_2.a_inv = "false";
defparam carry_12_1__ADD_2.PCK_LOCATION = "C18R4.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .PCK_LOCATION = "C20R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5]|qx_net  ),
	. di ( \ii2468|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[5] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t8_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_sc_vs_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.PCK_LOCATION = "C20R22.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t8_out1_reg.always_en = 1;
ADD1_A carry_12_1__ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3]|qx_net  ),
	. ci ( \carry_12_1__ADD_2|co_net  ),
	. co ( \carry_12_1__ADD_3|co_net  ),
	. s ( \carry_12_1__ADD_3|s_net  )
);
defparam carry_12_1__ADD_3.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_3.a_inv = "false";
defparam carry_12_1__ADD_3.PCK_LOCATION = "C18R4.lp0.add2.add0";
ADD1_A carry_12_1__ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4]|qx_net  ),
	. ci ( \carry_12_1__ADD_3|co_net  ),
	. co ( \carry_12_1__ADD_4|co_net  ),
	. s ( \carry_12_1__ADD_4|s_net  )
);
defparam carry_12_1__ADD_4.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_4.a_inv = "false";
defparam carry_12_1__ADD_4.PCK_LOCATION = "C18R4.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_4__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[25] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0]|qx_net  ),
	. di ( \ii2439|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[0] .always_en = 1;
ADD1_A carry_12_1__ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5]|qx_net  ),
	. ci ( \carry_12_1__ADD_4|co_net  ),
	. co ( \carry_12_1__ADD_5|co_net  ),
	. s ( \carry_12_1__ADD_5|s_net  )
);
defparam carry_12_1__ADD_5.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_5.a_inv = "false";
defparam carry_12_1__ADD_5.PCK_LOCATION = "C18R4.lp0.add2.add0";
ADD1_A carry_12_1__ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6]|qx_net  ),
	. ci ( \carry_12_1__ADD_5|co_net  ),
	. co ( \carry_12_1__ADD_6|co_net  ),
	. s ( \carry_12_1__ADD_6|s_net  )
);
defparam carry_12_1__ADD_6.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_6.a_inv = "false";
defparam carry_12_1__ADD_6.PCK_LOCATION = "C18R4.lp0.add2.add0";
REG mcu_arbiter_apb_sel_reg (
	. qx ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. di ( \ii3317|xy_net  ),
	. sr ( ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_apb_sel_reg.latch_mode = 0;
defparam mcu_arbiter_apb_sel_reg.init = 0;
defparam mcu_arbiter_apb_sel_reg.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_apb_sel_reg.sr_inv = 0;
defparam mcu_arbiter_apb_sel_reg.sync_mode = 1;
defparam mcu_arbiter_apb_sel_reg.no_sr = 1;
defparam mcu_arbiter_apb_sel_reg.sr_value = 0;
defparam mcu_arbiter_apb_sel_reg.PCK_LOCATION = "C4R20.lp0.reg0";
defparam mcu_arbiter_apb_sel_reg.clk_inv = 0;
defparam mcu_arbiter_apb_sel_reg.en_inv = 0;
defparam mcu_arbiter_apb_sel_reg.always_en = 1;
ADD1_A carry_12_1__ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7]|qx_net  ),
	. ci ( \carry_12_1__ADD_6|co_net  ),
	. co ( \carry_12_1__ADD_7|co_net  ),
	. s ( \carry_12_1__ADD_7|s_net  )
);
defparam carry_12_1__ADD_7.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_7.a_inv = "false";
defparam carry_12_1__ADD_7.PCK_LOCATION = "C18R4.lp0.add2.add0";
REG glue_rx_packet_tx_packet_fifo_sync_readen_reg (
	. qx ( \glue_rx_packet_tx_packet_fifo_sync_readen_reg|qx_net  ),
	. di ( \ii2140|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.init = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.PLACE_LOCATION = "C14R15.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.PCK_LOCATION = "C14R15.lp0.reg0";
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_readen_reg.always_en = 1;
ADD1_A carry_12_1__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8]|qx_net  ),
	. ci ( \carry_12_1__ADD_7|co_net  ),
	. co ( \carry_12_1__ADD_8|co_net  ),
	. s ( \carry_12_1__ADD_8|s_net  )
);
defparam carry_12_1__ADD_8.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_8.a_inv = "false";
defparam carry_12_1__ADD_8.PCK_LOCATION = "C18R5.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .PCK_LOCATION = "C10R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .PCK_LOCATION = "C20R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11] .always_en = 0;
ADD1_A carry_12_1__ADD_9 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9]|qx_net  ),
	. ci ( \carry_12_1__ADD_8|co_net  ),
	. co ( \carry_12_1__ADD_9|co_net  ),
	. s ( \carry_12_1__ADD_9|s_net  )
);
defparam carry_12_1__ADD_9.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_9.a_inv = "false";
defparam carry_12_1__ADD_9.PCK_LOCATION = "C18R5.lp0.add2.add0";
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc380 ,
		/* a_mac_out [23] (nc) */ nc381 ,
		/* a_mac_out [22] (nc) */ nc382 ,
		/* a_mac_out [21] (nc) */ nc383 ,
		/* a_mac_out [20] (nc) */ nc384 ,
		/* a_mac_out [19] (nc) */ nc385 ,
		/* a_mac_out [18] (nc) */ nc386 ,
		/* a_mac_out [17] (nc) */ nc387 ,
		/* a_mac_out [16] (nc) */ nc388 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc389 ,
		/* a_mac_out [2] (nc) */ nc390 ,
		/* a_mac_out [1] (nc) */ nc391 ,
		/* a_mac_out [0] (nc) */ nc392 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.PLACE_LOCATION = "C22R25.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.PCK_LOCATION = "C22R25.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0.amac_output_mode = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3]|qx_net  ),
	. di ( \ii3371|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6]|qx_net  ),
	. di ( \ii2469|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .PCK_LOCATION = "C6R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .PCK_LOCATION = "C20R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[26] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8]|qx_net  ),
	. di ( \ii3079|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In2p_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1]|qx_net  ),
	. di ( \ii2440|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[30] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .PCK_LOCATION = "C20R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12] .always_en = 0;
REG glue_rx_packet_tx_packet_u_scaler_t61_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t61_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.PLACE_LOCATION = "C20R26.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.PCK_LOCATION = "C20R26.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t61_out1_reg.always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[0]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[0]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[0] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4]|qx_net  ),
	. di ( \ii3384|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7]|qx_net  ),
	. di ( \ii2470|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .PCK_LOCATION = "C6R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_2_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .PCK_LOCATION = "C6R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .PLACE_LOCATION = "C14R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .PCK_LOCATION = "C14R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[27] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2]|qx_net  ),
	. di ( \ii2441|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[2] .always_en = 1;
REG glue_rd_start_f_reg (
	. qx ( \glue_rd_start_f_reg|qx_net  ),
	. di ( \ii2138|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rd_start_f_reg.latch_mode = 0;
defparam glue_rd_start_f_reg.init = 0;
defparam glue_rd_start_f_reg.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam glue_rd_start_f_reg.sr_inv = 1;
defparam glue_rd_start_f_reg.sync_mode = 0;
defparam glue_rd_start_f_reg.no_sr = 0;
defparam glue_rd_start_f_reg.sr_value = 0;
defparam glue_rd_start_f_reg.PCK_LOCATION = "C16R17.lp0.reg0";
defparam glue_rd_start_f_reg.clk_inv = 0;
defparam glue_rd_start_f_reg.en_inv = 0;
defparam glue_rd_start_f_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[31] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .PCK_LOCATION = "C20R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13] .always_en = 0;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg|qx_net  ),
	. di ( \ii2149|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.PCK_LOCATION = "C14R29.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg.always_en = 1;
LUT6 ii3195 (
	. xy ( \ii3195|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_8__ADD_8|co_net  )
);
defparam ii3195.PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.lut_0";
defparam ii3195.PCK_LOCATION = "C20R13.lp0.lut_0";
defparam ii3195.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[1]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[1]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[1] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5]|qx_net  ),
	. di ( \ii3385|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[6] .always_en = 1;
REG glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. di ( \ii3313|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.PCK_LOCATION = "C14R20.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .PCK_LOCATION = "C6R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3]|qx_net  ),
	. di ( \ii2442|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[3] .always_en = 1;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc393 ,
		/* a_mac_out [23] (nc) */ nc394 ,
		/* a_mac_out [22] (nc) */ nc395 ,
		/* a_mac_out [21] (nc) */ nc396 ,
		/* a_mac_out [20] (nc) */ nc397 ,
		/* a_mac_out [19] (nc) */ nc398 ,
		/* a_mac_out [18] (nc) */ nc399 ,
		/* a_mac_out [17] (nc) */ nc400 ,
		/* a_mac_out [16] (nc) */ nc401 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc402 ,
		/* a_mac_out [2] (nc) */ nc403 ,
		/* a_mac_out [1] (nc) */ nc404 ,
		/* a_mac_out [0] (nc) */ nc405 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.PLACE_LOCATION = "C22R15.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.PCK_LOCATION = "C22R15.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[3] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0]|qx_net  ),
	. di ( \ii2519|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[2]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[2]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[2] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6]|qx_net  ),
	. di ( \ii3371|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In3p_reg[7] .always_en = 1;
ADD1_A carry_9_12__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_12__ADD_0|co_net  ),
	. s ( \carry_9_12__ADD_0|s_net  )
);
defparam carry_9_12__ADD_0.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_0.a_inv = "true";
defparam carry_9_12__ADD_0.PCK_LOCATION = "C16R14.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .PCK_LOCATION = "C8R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .PCK_LOCATION = "C8R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[30] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t5_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.PCK_LOCATION = "C20R19.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t5_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4]|qx_net  ),
	. di ( \ii2443|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[4] .always_en = 1;
ADD1_A carry_9_12__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1]|qx_net  ),
	. ci ( \carry_9_12__ADD_0|co_net  ),
	. co ( \carry_9_12__ADD_1|co_net  ),
	. s ( \carry_9_12__ADD_1|s_net  )
);
defparam carry_9_12__ADD_1.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_1.a_inv = "true";
defparam carry_9_12__ADD_1.PCK_LOCATION = "C16R14.lp0.add2.add0";
ADD1_A carry_9_12__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2]|qx_net  ),
	. ci ( \carry_9_12__ADD_1|co_net  ),
	. co ( \carry_9_12__ADD_2|co_net  ),
	. s ( \carry_9_12__ADD_2|s_net  )
);
defparam carry_9_12__ADD_2.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_2.a_inv = "true";
defparam carry_9_12__ADD_2.PCK_LOCATION = "C16R14.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_9__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0] .always_en = 1;
ADD1_A carry_9_12__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3]|qx_net  ),
	. ci ( \carry_9_12__ADD_2|co_net  ),
	. co ( \carry_9_12__ADD_3|co_net  ),
	. s ( \carry_9_12__ADD_3|s_net  )
);
defparam carry_9_12__ADD_3.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_3.a_inv = "true";
defparam carry_9_12__ADD_3.PCK_LOCATION = "C16R14.lp0.add2.add0";
ADD1_A carry_9_12__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4]|qx_net  ),
	. ci ( \carry_9_12__ADD_3|co_net  ),
	. co ( \carry_9_12__ADD_4|co_net  ),
	. s ( \carry_9_12__ADD_4|s_net  )
);
defparam carry_9_12__ADD_4.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_4.a_inv = "true";
defparam carry_9_12__ADD_4.PCK_LOCATION = "C16R14.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[4] .always_en = 1;
LUT6 ii3224 (
	. xy ( \ii3224|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_9__ADD_8|co_net  )
);
defparam ii3224.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii3224.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii3224.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[3]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1]|qx_net  ),
	. di ( \ii2520|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1] .always_en = 1;
ADD1_A carry_9_12__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5]|qx_net  ),
	. ci ( \carry_9_12__ADD_4|co_net  ),
	. co ( \carry_9_12__ADD_5|co_net  ),
	. s ( \carry_9_12__ADD_5|s_net  )
);
defparam carry_9_12__ADD_5.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_5.a_inv = "true";
defparam carry_9_12__ADD_5.PCK_LOCATION = "C16R14.lp0.add2.add0";
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[3]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[3]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[3] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7] .always_en = 0;
ADD1_A carry_9_12__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6]|qx_net  ),
	. ci ( \carry_9_12__ADD_5|co_net  ),
	. co ( \carry_9_12__ADD_6|co_net  ),
	. s ( \carry_9_12__ADD_6|s_net  )
);
defparam carry_9_12__ADD_6.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_6.a_inv = "true";
defparam carry_9_12__ADD_6.PCK_LOCATION = "C16R14.lp0.add2.add0";
ADD1_A carry_9_12__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7]|qx_net  ),
	. ci ( \carry_9_12__ADD_6|co_net  ),
	. co ( \carry_9_12__ADD_7|co_net  ),
	. s ( \carry_9_12__ADD_7|s_net  )
);
defparam carry_9_12__ADD_7.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_7.a_inv = "true";
defparam carry_9_12__ADD_7.PCK_LOCATION = "C16R14.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t38_out1_reg[9] .always_en = 1;
ADD1_A carry_9_12__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_12__ADD_7|co_net  ),
	. co ( \carry_9_12__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_12__ADD_8.PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_12__ADD_8.a_inv = "false";
defparam carry_9_12__ADD_8.PCK_LOCATION = "C16R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .PCK_LOCATION = "C8R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t37_out1_reg[31] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[26]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5]|qx_net  ),
	. di ( \ii2444|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_9__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0]|qx_net  ),
	. di ( \ii2929|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .PCK_LOCATION = "C20R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .PCK_LOCATION = "C20R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In1p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2]|qx_net  ),
	. di ( \ii2521|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[4]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[4]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[4] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6]|qx_net  ),
	. di ( \ii2445|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[6] .always_en = 1;
REG glue_rx_packet_tx_packet_rstrf_reg (
	. qx ( \glue_rx_packet_tx_packet_rstrf_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_sc1_rstf_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rstrf_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.init = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rstrf_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rstrf_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.PCK_LOCATION = "C20R9.lp0.reg0";
defparam glue_rx_packet_tx_packet_rstrf_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rstrf_reg.always_en = 1;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc406 ,
		/* a_mac_out [23] (nc) */ nc407 ,
		/* a_mac_out [22] (nc) */ nc408 ,
		/* a_mac_out [21] (nc) */ nc409 ,
		/* a_mac_out [20] (nc) */ nc410 ,
		/* a_mac_out [19] (nc) */ nc411 ,
		/* a_mac_out [18] (nc) */ nc412 ,
		/* a_mac_out [17] (nc) */ nc413 ,
		/* a_mac_out [16] (nc) */ nc414 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc415 ,
		/* a_mac_out [2] (nc) */ nc416 ,
		/* a_mac_out [1] (nc) */ nc417 ,
		/* a_mac_out [0] (nc) */ nc418 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.PLACE_LOCATION = "C22R17.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.PCK_LOCATION = "C22R17.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_9__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1]|qx_net  ),
	. di ( \ii2930|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .PCK_LOCATION = "C20R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3]|qx_net  ),
	. di ( \ii2522|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[5]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[5]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[5] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7]|qx_net  ),
	. di ( \ii2446|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_11_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_9__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[3] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .PCK_LOCATION = "C4R6.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10] .always_en = 1;
LUT6 ii3253 (
	. xy ( \ii3253|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_10__ADD_8|co_net  )
);
defparam ii3253.PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.lut_0";
defparam ii3253.PCK_LOCATION = "C20R12.lp0.lut_0";
defparam ii3253.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2]|qx_net  ),
	. di ( \ii2931|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .PCK_LOCATION = "C20R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4]|qx_net  ),
	. di ( \ii2523|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4] .always_en = 1;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[16]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[6]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[6]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10]|qx_net  ),
	. di ( \ii2154|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_9__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[4] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11] .always_en = 1;
REG glue_pasm_packet_finish_reg (
	. qx ( \glue_pasm_packet_finish_reg|qx_net  ),
	. di ( \ii2135|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_pasm_packet_finish_reg.latch_mode = 0;
defparam glue_pasm_packet_finish_reg.init = 0;
defparam glue_pasm_packet_finish_reg.PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam glue_pasm_packet_finish_reg.sr_inv = 1;
defparam glue_pasm_packet_finish_reg.sync_mode = 0;
defparam glue_pasm_packet_finish_reg.no_sr = 0;
defparam glue_pasm_packet_finish_reg.sr_value = 0;
defparam glue_pasm_packet_finish_reg.PCK_LOCATION = "C10R22.lp0.reg0";
defparam glue_pasm_packet_finish_reg.clk_inv = 0;
defparam glue_pasm_packet_finish_reg.en_inv = 0;
defparam glue_pasm_packet_finish_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3]|qx_net  ),
	. di ( \ii2932|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .PCK_LOCATION = "C20R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5]|qx_net  ),
	. di ( \ii2524|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5] .always_en = 1;
ADD1_A carry_11_ADD_10 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \GND_0_inst|Y_net  ),
	. ci ( \carry_11_ADD_9|co_net  ),
	. co ( ),
	. s ( \carry_11_ADD_10|s_net  )
);
defparam carry_11_ADD_10.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_10.a_inv = "false";
defparam carry_11_ADD_10.PCK_LOCATION = "C18R18.lp0.add2.add0";
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[7]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[7]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memdatao_comb[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[7] .always_en = 0;
REG glue_rx_packet_tx_packet_u_data_process_first_3e_reg (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_first_3e_reg|qx_net  ),
	. di ( \ii2428|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.PCK_LOCATION = "C8R6.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_first_3e_reg.always_en = 1;
REG glue_rx_packet_tx_packet_tx_vsync_fo_reg (
	. qx ( \glue_rx_packet_tx_packet_tx_vsync_fo_reg|qx_net  ),
	. di ( \ii2424|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.init = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_tx_vsync_fo_reg.always_en = 1;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc419 ,
		/* a_mac_out [23] (nc) */ nc420 ,
		/* a_mac_out [22] (nc) */ nc421 ,
		/* a_mac_out [21] (nc) */ nc422 ,
		/* a_mac_out [20] (nc) */ nc423 ,
		/* a_mac_out [19] (nc) */ nc424 ,
		/* a_mac_out [18] (nc) */ nc425 ,
		/* a_mac_out [17] (nc) */ nc426 ,
		/* a_mac_out [16] (nc) */ nc427 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc428 ,
		/* a_mac_out [2] (nc) */ nc429 ,
		/* a_mac_out [1] (nc) */ nc430 ,
		/* a_mac_out [0] (nc) */ nc431 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.PLACE_LOCATION = "C22R11.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.PCK_LOCATION = "C22R11.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0.amac_output_mode = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10]|qx_net  ),
	. di ( \ii2409|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10] .always_en = 0;
REG \glue_cmd_s_reg[0]  (
	. qx ( \glue_cmd_s_reg[0]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[0] .latch_mode = 0;
defparam \glue_cmd_s_reg[0] .init = 0;
defparam \glue_cmd_s_reg[0] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[0] .sr_inv = 1;
defparam \glue_cmd_s_reg[0] .sync_mode = 0;
defparam \glue_cmd_s_reg[0] .no_sr = 0;
defparam \glue_cmd_s_reg[0] .sr_value = 0;
defparam \glue_cmd_s_reg[0] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_cmd_s_reg[0] .clk_inv = 0;
defparam \glue_cmd_s_reg[0] .en_inv = 0;
defparam \glue_cmd_s_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11]|qx_net  ),
	. di ( \ii2155|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11] .always_en = 0;
REG \glue_dnum_s_reg[10]  (
	. qx ( \glue_dnum_s_reg[10]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[18]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[10] .latch_mode = 0;
defparam \glue_dnum_s_reg[10] .init = 0;
defparam \glue_dnum_s_reg[10] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[10] .sr_inv = 1;
defparam \glue_dnum_s_reg[10] .sync_mode = 0;
defparam \glue_dnum_s_reg[10] .no_sr = 0;
defparam \glue_dnum_s_reg[10] .sr_value = 0;
defparam \glue_dnum_s_reg[10] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_dnum_s_reg[10] .clk_inv = 0;
defparam \glue_dnum_s_reg[10] .en_inv = 0;
defparam \glue_dnum_s_reg[10] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_9__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[5] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t85_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t85_out1_reg|qx_net  ),
	. di ( \ii2928|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.PLACE_LOCATION = "C6R23.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.PCK_LOCATION = "C6R23.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t85_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4]|qx_net  ),
	. di ( \ii2933|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .PCK_LOCATION = "C20R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6]|qx_net  ),
	. di ( \ii2525|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[8]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[8]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[8] .always_en = 0;
MIPI_PLL mipi_inst_u_mipi_pll (
	. CLKEXT ( ),
	. CLKREF ( \u_osc|OSC_net  ),
	. CM ( {
		/* CM [7] */ \mipi_inst_u_mipi2|CM[7]_net ,
		/* CM [6] */ \mipi_inst_u_mipi2|CM[6]_net ,
		/* CM [5] */ \mipi_inst_u_mipi2|CM[5]_net ,
		/* CM [4] */ \mipi_inst_u_mipi2|CM[4]_net ,
		/* CM [3] */ \mipi_inst_u_mipi2|CM[3]_net ,
		/* CM [2] */ \mipi_inst_u_mipi2|CM[2]_net ,
		/* CM [1] */ \mipi_inst_u_mipi2|CM[1]_net ,
		/* CM [0] */ \mipi_inst_u_mipi2|CM[0]_net 
	} ),
	. CN ( {
		/* CN [4] */ \mipi_inst_u_mipi2|CN[4]_net ,
		/* CN [3] */ \mipi_inst_u_mipi2|CN[3]_net ,
		/* CN [2] */ \mipi_inst_u_mipi2|CN[2]_net ,
		/* CN [1] */ \mipi_inst_u_mipi2|CN[1]_net ,
		/* CN [0] */ \mipi_inst_u_mipi2|CN[0]_net 
	} ),
	. CO ( {
		/* CO [1] */ \mipi_inst_u_mipi2|CO[1]_net ,
		/* CO [0] */ \mipi_inst_u_mipi2|CO[0]_net 
	} ),
	. PD_PLL ( \ii2049|xy_net  ),
	. CLKOUT1 ( \mipi_inst_u_mipi_pll|CLKOUT1_net  ),
	. CLKOUT2 ( \mipi_inst_u_mipi_pll|CLKOUT2_net  ),
	. LOCK ( \mipi_inst_u_mipi_pll|LOCK_net  )
);
defparam mipi_inst_u_mipi_pll.PLACE_LOCATION = "C2R8.mipi_wrap.mipi_pll";
defparam mipi_inst_u_mipi_pll.BYPASS_PLL = 0;
defparam mipi_inst_u_mipi_pll.PCK_LOCATION = "NONE";
defparam mipi_inst_u_mipi_pll.TST = 9;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[2] .always_en = 1;
GBUF u_gbuf_u_gbuf (
	. in ( \u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly|xy_net  ),
	. out ( \u_gbuf_u_gbuf|out_net  )
);
defparam u_gbuf_u_gbuf.PLACE_LOCATION = "NONE";
defparam u_gbuf_u_gbuf.M5_PRIM = "bool true";
defparam u_gbuf_u_gbuf.PCK_LOCATION = "NONE";
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11]|qx_net  ),
	. di ( \ii2410|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11] .always_en = 0;
REG glue_rx_packet_tx_packet_rx_payload_valid_d_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_valid_d_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload_valid_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.PCK_LOCATION = "C14R8.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_d_reg.always_en = 1;
REG \glue_cmd_s_reg[1]  (
	. qx ( \glue_cmd_s_reg[1]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[1] .latch_mode = 0;
defparam \glue_cmd_s_reg[1] .init = 0;
defparam \glue_cmd_s_reg[1] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[1] .sr_inv = 1;
defparam \glue_cmd_s_reg[1] .sync_mode = 0;
defparam \glue_cmd_s_reg[1] .no_sr = 0;
defparam \glue_cmd_s_reg[1] .sr_value = 0;
defparam \glue_cmd_s_reg[1] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_cmd_s_reg[1] .clk_inv = 0;
defparam \glue_cmd_s_reg[1] .en_inv = 0;
defparam \glue_cmd_s_reg[1] .always_en = 0;
REG mcu_arbiter_fifo_wr_d_reg (
	. qx ( \mcu_arbiter_fifo_wr_d_reg|qx_net  ),
	. di ( \ii3320|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_fifo_wr_d_reg.latch_mode = 0;
defparam mcu_arbiter_fifo_wr_d_reg.init = 0;
defparam mcu_arbiter_fifo_wr_d_reg.PLACE_LOCATION = "C6R18.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_fifo_wr_d_reg.sr_inv = 1;
defparam mcu_arbiter_fifo_wr_d_reg.sync_mode = 0;
defparam mcu_arbiter_fifo_wr_d_reg.no_sr = 0;
defparam mcu_arbiter_fifo_wr_d_reg.sr_value = 0;
defparam mcu_arbiter_fifo_wr_d_reg.PCK_LOCATION = "C6R18.lp0.reg0";
defparam mcu_arbiter_fifo_wr_d_reg.clk_inv = 0;
defparam mcu_arbiter_fifo_wr_d_reg.en_inv = 0;
defparam mcu_arbiter_fifo_wr_d_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12]|qx_net  ),
	. di ( \ii2156|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12] .always_en = 0;
REG \glue_dnum_s_reg[11]  (
	. qx ( \glue_dnum_s_reg[11]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[19]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[11] .latch_mode = 0;
defparam \glue_dnum_s_reg[11] .init = 0;
defparam \glue_dnum_s_reg[11] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[11] .sr_inv = 1;
defparam \glue_dnum_s_reg[11] .sync_mode = 0;
defparam \glue_dnum_s_reg[11] .no_sr = 0;
defparam \glue_dnum_s_reg[11] .sr_value = 0;
defparam \glue_dnum_s_reg[11] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_dnum_s_reg[11] .clk_inv = 0;
defparam \glue_dnum_s_reg[11] .en_inv = 0;
defparam \glue_dnum_s_reg[11] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_9__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[6] .always_en = 1;
LUT6 ii3282 (
	. xy ( \ii3282|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \carry_9_11__ADD_8|co_net  )
);
defparam ii3282.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii3282.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii3282.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13] .always_en = 1;
LUT6 ii3283 (
	. xy ( \ii3283|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_tx_vsync_fo_reg|qx_net  )
);
defparam ii3283.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3283.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3283.config_data = 64'b1010111010101110101011101010111010101110101011101010111010101110;
REG \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5]|qx_net  ),
	. di ( \ii2934|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .PCK_LOCATION = "C20R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[5] .always_en = 1;
LUT6 ii3284 (
	. xy ( \ii3284|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_tx_hsync_fo_reg|qx_net  )
);
defparam ii3284.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3284.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3284.config_data = 64'b1000100011111000100010001111100010001000111110001000100011111000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7]|qx_net  ),
	. di ( \ii2526|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7] .always_en = 1;
LUT6 ii3285 (
	. xy ( \ii3285|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0]|qx_net  )
);
defparam ii3285.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3285.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3285.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[9]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[9]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[3] .always_en = 1;
REG \glue_cmd_s_reg[2]  (
	. qx ( \glue_cmd_s_reg[2]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[2] .latch_mode = 0;
defparam \glue_cmd_s_reg[2] .init = 0;
defparam \glue_cmd_s_reg[2] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[2] .sr_inv = 1;
defparam \glue_cmd_s_reg[2] .sync_mode = 0;
defparam \glue_cmd_s_reg[2] .no_sr = 0;
defparam \glue_cmd_s_reg[2] .sr_value = 0;
defparam \glue_cmd_s_reg[2] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_cmd_s_reg[2] .clk_inv = 0;
defparam \glue_cmd_s_reg[2] .en_inv = 0;
defparam \glue_cmd_s_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13]|qx_net  ),
	. di ( \ii2157|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13] .always_en = 0;
REG \glue_dnum_s_reg[12]  (
	. qx ( \glue_dnum_s_reg[12]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[20]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[12] .latch_mode = 0;
defparam \glue_dnum_s_reg[12] .init = 0;
defparam \glue_dnum_s_reg[12] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[12] .sr_inv = 1;
defparam \glue_dnum_s_reg[12] .sync_mode = 0;
defparam \glue_dnum_s_reg[12] .no_sr = 0;
defparam \glue_dnum_s_reg[12] .sr_value = 0;
defparam \glue_dnum_s_reg[12] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_dnum_s_reg[12] .clk_inv = 0;
defparam \glue_dnum_s_reg[12] .en_inv = 0;
defparam \glue_dnum_s_reg[12] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_9__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[7] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[10]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[10]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[10] .always_en = 1;
REG glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. di ( \ii3316|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.PCK_LOCATION = "C14R20.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg.always_en = 1;
LUT6 ii3304 (
	. xy ( \ii3304|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_1|s_net  )
);
defparam ii3304.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3304.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3304.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .PLACE_LOCATION = "C8R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .PCK_LOCATION = "C8R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0] .always_en = 1;
LUT6 ii3305 (
	. xy ( \ii3305|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_2|s_net  )
);
defparam ii3305.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3305.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3305.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
H6_MAC glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0 (
	. a_acc_en ( \GND_0_inst|Y_net  ),
	. a_dinx ( {
		/* a_dinx [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net ,
		/* a_dinx [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net ,
		/* a_dinx [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net ,
		/* a_dinx [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net ,
		/* a_dinx [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net ,
		/* a_dinx [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net ,
		/* a_dinx [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7]|qx_net ,
		/* a_dinx [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6]|qx_net ,
		/* a_dinx [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5]|qx_net ,
		/* a_dinx [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4]|qx_net ,
		/* a_dinx [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3]|qx_net ,
		/* a_dinx [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2]|qx_net ,
		/* a_dinx [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1]|qx_net ,
		/* a_dinx [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0]|qx_net 
	} ),
	. a_dinxy_cen ( \VCC_0_inst|Y_net  ),
	. a_diny ( {
		/* a_diny [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net ,
		/* a_diny [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net ,
		/* a_diny [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net ,
		/* a_diny [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net ,
		/* a_diny [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[5]|qx_net ,
		/* a_diny [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[4]|qx_net ,
		/* a_diny [3] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3]|qx_net ,
		/* a_diny [2] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2]|qx_net ,
		/* a_diny [1] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1]|qx_net ,
		/* a_diny [0] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0]|qx_net 
	} ),
	. a_dinz ( {
		/* a_dinz [24] */ \GND_0_inst|Y_net ,
		/* a_dinz [23] */ \GND_0_inst|Y_net ,
		/* a_dinz [22] */ \GND_0_inst|Y_net ,
		/* a_dinz [21] */ \GND_0_inst|Y_net ,
		/* a_dinz [20] */ \GND_0_inst|Y_net ,
		/* a_dinz [19] */ \GND_0_inst|Y_net ,
		/* a_dinz [18] */ \GND_0_inst|Y_net ,
		/* a_dinz [17] */ \GND_0_inst|Y_net ,
		/* a_dinz [16] */ \GND_0_inst|Y_net ,
		/* a_dinz [15] */ \GND_0_inst|Y_net ,
		/* a_dinz [14] */ \GND_0_inst|Y_net ,
		/* a_dinz [13] */ \GND_0_inst|Y_net ,
		/* a_dinz [12] */ \GND_0_inst|Y_net ,
		/* a_dinz [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7]|qx_net ,
		/* a_dinz [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6]|qx_net ,
		/* a_dinz [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5]|qx_net ,
		/* a_dinz [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4]|qx_net ,
		/* a_dinz [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3]|qx_net ,
		/* a_dinz [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2]|qx_net ,
		/* a_dinz [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1]|qx_net ,
		/* a_dinz [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0]|qx_net ,
		/* a_dinz [3] */ \GND_0_inst|Y_net ,
		/* a_dinz [2] */ \GND_0_inst|Y_net ,
		/* a_dinz [1] */ \GND_0_inst|Y_net ,
		/* a_dinz [0] */ \GND_0_inst|Y_net 
	} ),
	. a_dinz_cen ( \VCC_0_inst|Y_net  ),
	. a_dinz_en ( \VCC_0_inst|Y_net  ),
	. a_in_sr ( \VCC_0_inst|Y_net  ),
	. a_mac_out_cen ( \VCC_0_inst|Y_net  ),
	. a_out_sr ( \VCC_0_inst|Y_net  ),
	. a_sload ( \GND_0_inst|Y_net  ),
	. b_acc_en ( ),
	. b_dinx ( )
,
	. b_dinxy_cen ( ),
	. b_diny ( )
,
	. b_dinz ( )
,
	. b_dinz_cen ( ),
	. b_dinz_en ( ),
	. b_in_sr ( ),
	. b_mac_out_cen ( ),
	. b_out_sr ( ),
	. b_sload ( ),
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. dsp_en ( ),
	. a_mac_out ( {
		/* a_mac_out [24] (nc) */ nc432 ,
		/* a_mac_out [23] (nc) */ nc433 ,
		/* a_mac_out [22] (nc) */ nc434 ,
		/* a_mac_out [21] (nc) */ nc435 ,
		/* a_mac_out [20] (nc) */ nc436 ,
		/* a_mac_out [19] (nc) */ nc437 ,
		/* a_mac_out [18] (nc) */ nc438 ,
		/* a_mac_out [17] (nc) */ nc439 ,
		/* a_mac_out [16] (nc) */ nc440 ,
		/* a_mac_out [15] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net ,
		/* a_mac_out [14] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net ,
		/* a_mac_out [13] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net ,
		/* a_mac_out [12] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net ,
		/* a_mac_out [11] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[11]_net ,
		/* a_mac_out [10] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[10]_net ,
		/* a_mac_out [9] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[9]_net ,
		/* a_mac_out [8] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[8]_net ,
		/* a_mac_out [7] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[7]_net ,
		/* a_mac_out [6] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[6]_net ,
		/* a_mac_out [5] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[5]_net ,
		/* a_mac_out [4] */ \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[4]_net ,
		/* a_mac_out [3] (nc) */ nc441 ,
		/* a_mac_out [2] (nc) */ nc442 ,
		/* a_mac_out [1] (nc) */ nc443 ,
		/* a_mac_out [0] (nc) */ nc444 
	} ),
	. a_overflow ( ),
	. b_mac_out ( )
,
	. b_overflow ( )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.adiny_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.bdinx_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.a_out_rstn_sel = 48'b111111111111111111111111111111111111111111111111;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.a_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.bdinz_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.a_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.b_in_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.a_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.b_out_setn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.adinx_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.bmac_output_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.a_in_rstn_sel = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.b_in_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.modea_sel = 2;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.adinz_input_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.bdiny_input_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.b_out_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.b_sr_syn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.modeb_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.a_out_setn_sel = 48'b000000000000000000000000000000000000000000000000;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.PLACE_LOCATION = "C22R13.mac_guts.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.b_ovf_rstn_sel = 0;
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.PCK_LOCATION = "C22R13.mac";
defparam glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0.amac_output_mode = 0;
LUT6 ii3306 (
	. xy ( \ii3306|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_3|s_net  )
);
defparam ii3306.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3306.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3306.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii3307 (
	. xy ( \ii3307|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_4|s_net  )
);
defparam ii3307.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3307.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3307.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii3308 (
	. xy ( \ii3308|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_5|s_net  )
);
defparam ii3308.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3308.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3308.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[4] .always_en = 1;
LUT6 ii3309 (
	. xy ( \ii3309|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_6|s_net  )
);
defparam ii3309.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3309.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3309.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii3310 (
	. xy ( \ii3310|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \carry_8_ADD_7|s_net  )
);
defparam ii3310.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3310.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3310.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ),
	. di ( \ii2568|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .PCK_LOCATION = "C18R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0] .always_en = 1;
REG \glue_cmd_s_reg[3]  (
	. qx ( \glue_cmd_s_reg[3]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[3] .latch_mode = 0;
defparam \glue_cmd_s_reg[3] .init = 0;
defparam \glue_cmd_s_reg[3] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[3] .sr_inv = 1;
defparam \glue_cmd_s_reg[3] .sync_mode = 0;
defparam \glue_cmd_s_reg[3] .no_sr = 0;
defparam \glue_cmd_s_reg[3] .sr_value = 0;
defparam \glue_cmd_s_reg[3] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_cmd_s_reg[3] .clk_inv = 0;
defparam \glue_cmd_s_reg[3] .en_inv = 0;
defparam \glue_cmd_s_reg[3] .always_en = 0;
LUT6 ii3311 (
	. xy ( \ii3311|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0]|qx_net  )
);
defparam ii3311.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3311.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3311.config_data = 64'b0000000000000100000000000000000000000000000000000000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14]|qx_net  ),
	. di ( \ii2158|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14] .always_en = 0;
REG \glue_dnum_s_reg[13]  (
	. qx ( \glue_dnum_s_reg[13]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[21]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[13] .latch_mode = 0;
defparam \glue_dnum_s_reg[13] .init = 0;
defparam \glue_dnum_s_reg[13] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[13] .sr_inv = 1;
defparam \glue_dnum_s_reg[13] .sync_mode = 0;
defparam \glue_dnum_s_reg[13] .no_sr = 0;
defparam \glue_dnum_s_reg[13] .sr_value = 0;
defparam \glue_dnum_s_reg[13] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_dnum_s_reg[13] .clk_inv = 0;
defparam \glue_dnum_s_reg[13] .en_inv = 0;
defparam \glue_dnum_s_reg[13] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8]|qx_net  ),
	. di ( \ii3224|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .PCK_LOCATION = "C20R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In2p_reg[8] .always_en = 1;
LUT6 ii3312 (
	. xy ( \ii3312|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_tx_vsync_fo_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_tx_hsync_fo_reg|qx_net  ),
	. f0 ( \ii3311|xy_net  )
);
defparam ii3312.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3312.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3312.config_data = 64'b1111111111111111111111111111110111111100111111001111110011111100;
REG \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15]  (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .init = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15] .always_en = 1;
LUT6 ii3313 (
	. xy ( \ii3313|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_d_reg|qx_net  )
);
defparam ii3313.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3313.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3313.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[11]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[11]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[11] .always_en = 1;
LUT6 ii3314 (
	. xy ( \ii3314|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_tx_hsync_fo_reg|qx_net  )
);
defparam ii3314.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3314.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3314.config_data = 64'b1000100011111000100010001111100010001000111110001000100011111000;
REG \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1] .always_en = 1;
LUT6 ii3315 (
	. xy ( \ii3315|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_tx_hsync_fo_reg|qx_net  )
);
defparam ii3315.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3315.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3315.config_data = 64'b1000100011111000100010001111100010001000111110001000100011111000;
REG \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0]|qx_net  ),
	. di ( \ii3387|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0] .always_en = 0;
LUT6 ii3316 (
	. xy ( \ii3316|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg|qx_net  ),
	. f0 ( \ii3313|xy_net  )
);
defparam ii3316.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii3316.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii3316.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .PLACE_LOCATION = "C10R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .PCK_LOCATION = "C10R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0] .always_en = 1;
LUT6 ii3317 (
	. xy ( \ii3317|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[17]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[11]_net  )
);
defparam ii3317.PLACE_LOCATION = "C8R17.le_tile.le_guts.lp0.lut_0";
defparam ii3317.PCK_LOCATION = "C8R17.lp0.lut_0";
defparam ii3317.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0] .always_en = 1;
LUT6 ii3318 (
	. xy ( \ii3318|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|mempswr_comb_net  ),
	. f0 ( \u_8051_u_h6_8051|mempsrd_comb_net  )
);
defparam ii3318.PLACE_LOCATION = "C4R17.le_tile.le_guts.lp0.lut_0";
defparam ii3318.PCK_LOCATION = "C4R17.lp0.lut_0";
defparam ii3318.config_data = 64'b1110111011101110111011101110111011101110111011101110111011101110;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0]|qx_net  ),
	. di ( \ii2340|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .PCK_LOCATION = "C16R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[5] .always_en = 1;
LUT6 ii3319 (
	. xy ( \ii3319|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memwr_comb_net  ),
	. f0 ( \u_8051_u_h6_8051|memrd_comb_net  )
);
defparam ii3319.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.lut_0";
defparam ii3319.PCK_LOCATION = "C4R18.lp0.lut_0";
defparam ii3319.config_data = 64'b1110111011101110111011101110111011101110111011101110111011101110;
LUT6 ii3320 (
	. xy ( \ii3320|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f0 ( \ii2039|xy_net  )
);
defparam ii3320.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3320.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3320.config_data = 64'b0000001000000010000000100000001000000010000000100000001000000010;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1]|qx_net  ),
	. di ( \ii2569|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1] .always_en = 1;
REG \glue_cmd_s_reg[4]  (
	. qx ( \glue_cmd_s_reg[4]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[4] .latch_mode = 0;
defparam \glue_cmd_s_reg[4] .init = 0;
defparam \glue_cmd_s_reg[4] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[4] .sr_inv = 1;
defparam \glue_cmd_s_reg[4] .sync_mode = 0;
defparam \glue_cmd_s_reg[4] .no_sr = 0;
defparam \glue_cmd_s_reg[4] .sr_value = 0;
defparam \glue_cmd_s_reg[4] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_cmd_s_reg[4] .clk_inv = 0;
defparam \glue_cmd_s_reg[4] .en_inv = 0;
defparam \glue_cmd_s_reg[4] .always_en = 0;
LUT6 ii3321 (
	. xy ( \ii3321|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f0 ( \ii2039|xy_net  )
);
defparam ii3321.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii3321.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii3321.config_data = 64'b1000000010000000100000001000000010000000100000001000000010000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15]|qx_net  ),
	. di ( \ii2159|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15] .always_en = 0;
FIFO5K glue_rx_packet_tx_packet_fifo_sync_inst_u_inst (
	. dout ( {
		/* dout [15] (nc) */ nc445 ,
		/* dout [14] (nc) */ nc446 ,
		/* dout [13] (nc) */ nc447 ,
		/* dout [12] (nc) */ nc448 ,
		/* dout [11] (nc) */ nc449 ,
		/* dout [10] (nc) */ nc450 ,
		/* dout [9] (nc) */ nc451 ,
		/* dout [8] (nc) */ nc452 ,
		/* dout [7] (nc) */ nc453 ,
		/* dout [6] (nc) */ nc454 ,
		/* dout [5] (nc) */ nc455 ,
		/* dout [4] (nc) */ nc456 ,
		/* dout [3] (nc) */ nc457 ,
		/* dout [2] (nc) */ nc458 ,
		/* dout [1] */ \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|dout[1]_net ,
		/* dout [0] */ \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|dout[0]_net 
	} ),
	. doutp ( )
,
	. din ( {
		/* din [15] */ \GND_0_inst|Y_net ,
		/* din [14] */ \GND_0_inst|Y_net ,
		/* din [13] */ \GND_0_inst|Y_net ,
		/* din [12] */ \GND_0_inst|Y_net ,
		/* din [11] */ \GND_0_inst|Y_net ,
		/* din [10] */ \GND_0_inst|Y_net ,
		/* din [9] */ \GND_0_inst|Y_net ,
		/* din [8] */ \GND_0_inst|Y_net ,
		/* din [7] */ \GND_0_inst|Y_net ,
		/* din [6] */ \GND_0_inst|Y_net ,
		/* din [5] */ \GND_0_inst|Y_net ,
		/* din [4] */ \GND_0_inst|Y_net ,
		/* din [3] */ \GND_0_inst|Y_net ,
		/* din [2] */ \GND_0_inst|Y_net ,
		/* din [1] */ \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net ,
		/* din [0] */ \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net 
	} ),
	. dinp ( )
,
	. writeclk ( \u_pll_pll_u0|CO0_net  ),
	. readclk ( \u_gbuf_u_gbuf|out_net  ),
	. writeen ( \ii1983|xy_net  ),
	. readen ( \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|empty_net  ),
	. reset ( \ii1982_dup|xy_net  ),
	. regce ( ),
	. writesave ( \GND_0_inst|Y_net  ),
	. writedrop ( \GND_0_inst|Y_net  ),
	. full ( ),
	. empty ( \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|empty_net  ),
	. almostfull ( ),
	. almostempty ( ),
	. overflow ( ),
	. underflow ( ),
	. writedropflag ( )
);
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.readwidth = 4;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.PLACE_LOCATION = "C12R1.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core.bram5k_0";
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.writeclk_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.peek = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.PCK_LOCATION = "C12R1.u0_emb_top.emb18k_wrapper.u0_emb18k_core.bram5k_0";
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.readclk_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.outreg = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.writewidth = 4;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.almostfullth = 0;
defparam glue_rx_packet_tx_packet_fifo_sync_inst_u_inst.almostemptyth = 0;
REG \glue_dnum_s_reg[14]  (
	. qx ( \glue_dnum_s_reg[14]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[22]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[14] .latch_mode = 0;
defparam \glue_dnum_s_reg[14] .init = 0;
defparam \glue_dnum_s_reg[14] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[14] .sr_inv = 1;
defparam \glue_dnum_s_reg[14] .sync_mode = 0;
defparam \glue_dnum_s_reg[14] .no_sr = 0;
defparam \glue_dnum_s_reg[14] .sr_value = 0;
defparam \glue_dnum_s_reg[14] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_dnum_s_reg[14] .clk_inv = 0;
defparam \glue_dnum_s_reg[14] .en_inv = 0;
defparam \glue_dnum_s_reg[14] .always_en = 0;
LUT6 ii3322 (
	. xy ( \ii3322|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_mipi_sel_reg|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memdatao_comb[0]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f0 ( \ii2039|xy_net  )
);
defparam ii3322.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii3322.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii3322.config_data = 64'b1111111111011111001000000000000011111111110111110010000000000000;
REG mcu_arbiter_reg_memack_reg (
	. qx ( \mcu_arbiter_reg_memack_reg|qx_net  ),
	. di ( \ii3332|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_reg_memack_reg.latch_mode = 0;
defparam mcu_arbiter_reg_memack_reg.init = 0;
defparam mcu_arbiter_reg_memack_reg.PLACE_LOCATION = "C4R19.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_reg_memack_reg.sr_inv = 1;
defparam mcu_arbiter_reg_memack_reg.sync_mode = 0;
defparam mcu_arbiter_reg_memack_reg.no_sr = 0;
defparam mcu_arbiter_reg_memack_reg.sr_value = 0;
defparam mcu_arbiter_reg_memack_reg.PCK_LOCATION = "C4R19.lp0.reg0";
defparam mcu_arbiter_reg_memack_reg.clk_inv = 0;
defparam mcu_arbiter_reg_memack_reg.en_inv = 0;
defparam mcu_arbiter_reg_memack_reg.always_en = 1;
LUT6 ii3323 (
	. xy ( \ii3323|xy_net  ),
	. f5 ( \mcu_arbiter_mipi_sel_reg|qx_net  ),
	. f4 ( \mcu_arbiter_func_reg[0]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3323.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii3323.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii3323.config_data = 64'b0000000000110000000000000001000000000000001000000000000000000000;
REG mcu_arbiter_u_emif2apb_fpga_HRD_reg (
	. qx ( \mcu_arbiter_u_emif2apb_fpga_HRD_reg|qx_net  ),
	. di ( \ii3335|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.latch_mode = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.init = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.sr_inv = 1;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.sync_mode = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.no_sr = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.sr_value = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.PCK_LOCATION = "C4R16.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.clk_inv = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.en_inv = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HRD_reg.always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[12]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[12]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[12] .always_en = 1;
LUT6 ii3324 (
	. xy ( \ii3324|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memrd_comb_net  ),
	. f0 ( \ii2038|xy_net  )
);
defparam ii3324.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.lut_0";
defparam ii3324.PCK_LOCATION = "C4R18.lp0.lut_0";
defparam ii3324.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .PLACE_LOCATION = "C6R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .PCK_LOCATION = "C6R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2] .always_en = 1;
LUT6 ii3325 (
	. xy ( \ii3325|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[1]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3325.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.lut_0";
defparam ii3325.PCK_LOCATION = "C4R16.lp0.lut_0";
defparam ii3325.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
REG \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1] .always_en = 0;
LUT6 ii3326 (
	. xy ( \ii3326|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[2]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3326.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3326.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3326.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .PLACE_LOCATION = "C10R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .PCK_LOCATION = "C10R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1] .always_en = 1;
LUT6 ii3327 (
	. xy ( \ii3327|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[3]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3327.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3327.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3327.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1] .always_en = 1;
LUT6 ii3328 (
	. xy ( \ii3328|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[4]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3328.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3328.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3328.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1]|qx_net  ),
	. di ( \ii2370|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .PCK_LOCATION = "C16R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[1] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0]|qx_net  ),
	. di ( \ii2220|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[6] .always_en = 1;
LUT6 ii3329 (
	. xy ( \ii3329|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[5]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3329.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3329.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3329.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
LUT6 ii3330 (
	. xy ( \ii3330|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[6]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3330.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3330.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3330.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2]|qx_net  ),
	. di ( \ii2570|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2] .always_en = 1;
REG \glue_cmd_s_reg[5]  (
	. qx ( \glue_cmd_s_reg[5]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[5] .latch_mode = 0;
defparam \glue_cmd_s_reg[5] .init = 0;
defparam \glue_cmd_s_reg[5] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[5] .sr_inv = 1;
defparam \glue_cmd_s_reg[5] .sync_mode = 0;
defparam \glue_cmd_s_reg[5] .no_sr = 0;
defparam \glue_cmd_s_reg[5] .sr_value = 0;
defparam \glue_cmd_s_reg[5] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_cmd_s_reg[5] .clk_inv = 0;
defparam \glue_cmd_s_reg[5] .en_inv = 0;
defparam \glue_cmd_s_reg[5] .always_en = 0;
LUT6 ii3331 (
	. xy ( \ii3331|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_func_reg[7]|qx_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3331.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3331.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3331.config_data = 64'b0000000000100000000000000000000000000000001000000000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16]|qx_net  ),
	. di ( \ii2161|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16] .always_en = 0;
REG \glue_dnum_s_reg[15]  (
	. qx ( \glue_dnum_s_reg[15]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[23]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_dnum_s_reg[15] .latch_mode = 0;
defparam \glue_dnum_s_reg[15] .init = 0;
defparam \glue_dnum_s_reg[15] .PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.reg0";
defparam \glue_dnum_s_reg[15] .sr_inv = 1;
defparam \glue_dnum_s_reg[15] .sync_mode = 0;
defparam \glue_dnum_s_reg[15] .no_sr = 0;
defparam \glue_dnum_s_reg[15] .sr_value = 0;
defparam \glue_dnum_s_reg[15] .PCK_LOCATION = "C14R26.lp0.reg0";
defparam \glue_dnum_s_reg[15] .clk_inv = 0;
defparam \glue_dnum_s_reg[15] .en_inv = 0;
defparam \glue_dnum_s_reg[15] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .PCK_LOCATION = "C14R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[0] .always_en = 1;
LUT6 ii3332 (
	. xy ( \ii3332|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \ii3319|xy_net  ),
	. f0 ( \ii2038|xy_net  )
);
defparam ii3332.PLACE_LOCATION = "C4R19.le_tile.le_guts.lp0.lut_0";
defparam ii3332.PCK_LOCATION = "C4R19.lp0.lut_0";
defparam ii3332.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii3333 (
	. xy ( \ii3333|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memrd_comb_net  ),
	. f0 ( \ii3317|xy_net  )
);
defparam ii3333.PLACE_LOCATION = "C8R17.le_tile.le_guts.lp0.lut_0";
defparam ii3333.PCK_LOCATION = "C8R17.lp0.lut_0";
defparam ii3333.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[13]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[13]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[13] .always_en = 1;
ADD1_A carry_9_9__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_9__ADD_0|co_net  ),
	. s ( \carry_9_9__ADD_0|s_net  )
);
defparam carry_9_9__ADD_0.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_0.a_inv = "true";
defparam carry_9_9__ADD_0.PCK_LOCATION = "C18R13.lp0.add2.add0";
LUT6 ii3334 (
	. xy ( \ii3334|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mipi_inst_u_mipi2|pready_net  ),
	. f0 ( \mipi_inst_u_mipi1|pready_net  )
);
defparam ii3334.PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.lut_0";
defparam ii3334.PCK_LOCATION = "C4R15.lp0.lut_0";
defparam ii3334.config_data = 64'b1110111011101110111011101110111011101110111011101110111011101110;
ADD1_A carry_12_0__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_12_0__ADD_0|co_net  ),
	. s ( )
);
defparam carry_12_0__ADD_0.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_0.a_inv = "false";
defparam carry_12_0__ADD_0.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1]|qx_net  ),
	. ci ( \carry_9_9__ADD_0|co_net  ),
	. co ( \carry_9_9__ADD_1|co_net  ),
	. s ( \carry_9_9__ADD_1|s_net  )
);
defparam carry_9_9__ADD_1.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_1.a_inv = "true";
defparam carry_9_9__ADD_1.PCK_LOCATION = "C18R13.lp0.add2.add0";
LUT6 ii3335 (
	. xy ( \ii3335|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memrd_s_reg|qx_net  ),
	. f3 ( \mcu_arbiter_u_emif2apb_memack_reg|qx_net  ),
	. f2 ( \mcu_arbiter_u_emif2apb_fpga_HRD_reg|qx_net  ),
	. f1 ( \ii3334|xy_net  ),
	. f0 ( \ii3333|xy_net  )
);
defparam ii3335.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.lut_0";
defparam ii3335.PCK_LOCATION = "C4R16.lp0.lut_0";
defparam ii3335.config_data = 64'b0011000000110000001100000011001000110000001100000011000000110010;
REG \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2]|qx_net  ),
	. di ( \ii3386|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2] .always_en = 0;
ADD1_A carry_12_0__ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1]|qx_net  ),
	. ci ( \carry_12_0__ADD_0|co_net  ),
	. co ( \carry_12_0__ADD_1|co_net  ),
	. s ( \carry_12_0__ADD_1|s_net  )
);
defparam carry_12_0__ADD_1.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_1.a_inv = "false";
defparam carry_12_0__ADD_1.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2]|qx_net  ),
	. ci ( \carry_9_9__ADD_1|co_net  ),
	. co ( \carry_9_9__ADD_2|co_net  ),
	. s ( \carry_9_9__ADD_2|s_net  )
);
defparam carry_9_9__ADD_2.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_2.a_inv = "true";
defparam carry_9_9__ADD_2.PCK_LOCATION = "C18R13.lp0.add2.add0";
LUT6 ii3336 (
	. xy ( \ii3336|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \mcu_arbiter_u_emif2apb_memwr_s_reg|qx_net  ),
	. f2 ( \mcu_arbiter_u_emif2apb_memack_reg|qx_net  ),
	. f1 ( \u_8051_u_h6_8051|memwr_comb_net  ),
	. f0 ( \ii3317|xy_net  )
);
defparam ii3336.PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.lut_0";
defparam ii3336.PCK_LOCATION = "C4R15.lp0.lut_0";
defparam ii3336.config_data = 64'b0000000000001000000000000000100000000000000010000000000000001000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2] .always_en = 1;
ADD1_A carry_12_0__ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2]|qx_net  ),
	. ci ( \carry_12_0__ADD_1|co_net  ),
	. co ( \carry_12_0__ADD_2|co_net  ),
	. s ( \carry_12_0__ADD_2|s_net  )
);
defparam carry_12_0__ADD_2.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_2.a_inv = "false";
defparam carry_12_0__ADD_2.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3]|qx_net  ),
	. ci ( \carry_9_9__ADD_2|co_net  ),
	. co ( \carry_9_9__ADD_3|co_net  ),
	. s ( \carry_9_9__ADD_3|s_net  )
);
defparam carry_9_9__ADD_3.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_3.a_inv = "true";
defparam carry_9_9__ADD_3.PCK_LOCATION = "C18R13.lp0.add2.add0";
LUT6 ii3337 (
	. xy ( \ii3337|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1]|qx_net  ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0]|qx_net  )
);
defparam ii3337.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.lut_0";
defparam ii3337.PCK_LOCATION = "C4R16.lp0.lut_0";
defparam ii3337.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2] .always_en = 1;
ADD1_A carry_12_0__ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3]|qx_net  ),
	. ci ( \carry_12_0__ADD_2|co_net  ),
	. co ( \carry_12_0__ADD_3|co_net  ),
	. s ( \carry_12_0__ADD_3|s_net  )
);
defparam carry_12_0__ADD_3.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_3.a_inv = "false";
defparam carry_12_0__ADD_3.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4]|qx_net  ),
	. ci ( \carry_9_9__ADD_3|co_net  ),
	. co ( \carry_9_9__ADD_4|co_net  ),
	. s ( \carry_9_9__ADD_4|s_net  )
);
defparam carry_9_9__ADD_4.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_4.a_inv = "true";
defparam carry_9_9__ADD_4.PCK_LOCATION = "C18R13.lp0.add2.add0";
LUT6 ii3338 (
	. xy ( \ii3338|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg|qx_net  ),
	. f2 ( \ii3337|xy_net  ),
	. f1 ( \ii3334|xy_net  ),
	. f0 ( \ii3336|xy_net  )
);
defparam ii3338.PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.lut_0";
defparam ii3338.PCK_LOCATION = "C4R15.lp0.lut_0";
defparam ii3338.config_data = 64'b0011001100100000001100110010000000110011001000000011001100100000;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2]|qx_net  ),
	. di ( \ii2371|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .PCK_LOCATION = "C16R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1]|qx_net  ),
	. di ( \ii2231|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1] .always_en = 0;
ADD1_A carry_12_0__ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4]|qx_net  ),
	. ci ( \carry_12_0__ADD_3|co_net  ),
	. co ( \carry_12_0__ADD_4|co_net  ),
	. s ( \carry_12_0__ADD_4|s_net  )
);
defparam carry_12_0__ADD_4.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_4.a_inv = "false";
defparam carry_12_0__ADD_4.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5]|qx_net  ),
	. ci ( \carry_9_9__ADD_4|co_net  ),
	. co ( \carry_9_9__ADD_5|co_net  ),
	. s ( \carry_9_9__ADD_5|s_net  )
);
defparam carry_9_9__ADD_5.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_5.a_inv = "true";
defparam carry_9_9__ADD_5.PCK_LOCATION = "C18R13.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In3p_reg[7] .always_en = 1;
LUT6 ii3339 (
	. xy ( \ii3339|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg|qx_net  ),
	. f0 ( \ii3334|xy_net  )
);
defparam ii3339.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3339.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3339.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii3340 (
	. xy ( \ii3340|xy_net  ),
	. f5 ( \mcu_arbiter_u_emif2apb_memack_reg|qx_net  ),
	. f4 ( \ii3337|xy_net  ),
	. f3 ( \ii3319|xy_net  ),
	. f2 ( \ii3317|xy_net  ),
	. f1 ( \ii3339|xy_net  ),
	. f0 ( \ii3336|xy_net  )
);
defparam ii3340.PLACE_LOCATION = "C6R17.le_tile.le_guts.lp0.lut_0";
defparam ii3340.PCK_LOCATION = "C6R17.lp0.lut_0";
defparam ii3340.config_data = 64'b1111000000000000111100000000000011000000000000001110000000000000;
REG \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0]|qx_net  ),
	. di ( \ii3367|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3]|qx_net  ),
	. di ( \ii2571|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0]|qx_net  ),
	. di ( \ii2431|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .PCK_LOCATION = "C14R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0] .always_en = 1;
REG \glue_cmd_s_reg[6]  (
	. qx ( \glue_cmd_s_reg[6]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[6] .latch_mode = 0;
defparam \glue_cmd_s_reg[6] .init = 0;
defparam \glue_cmd_s_reg[6] .PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[6] .sr_inv = 1;
defparam \glue_cmd_s_reg[6] .sync_mode = 0;
defparam \glue_cmd_s_reg[6] .no_sr = 0;
defparam \glue_cmd_s_reg[6] .sr_value = 0;
defparam \glue_cmd_s_reg[6] .PCK_LOCATION = "C14R29.lp0.reg0";
defparam \glue_cmd_s_reg[6] .clk_inv = 0;
defparam \glue_cmd_s_reg[6] .en_inv = 0;
defparam \glue_cmd_s_reg[6] .always_en = 0;
ADD1_A carry_12_0__ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5]|qx_net  ),
	. ci ( \carry_12_0__ADD_4|co_net  ),
	. co ( \carry_12_0__ADD_5|co_net  ),
	. s ( \carry_12_0__ADD_5|s_net  )
);
defparam carry_12_0__ADD_5.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_5.a_inv = "false";
defparam carry_12_0__ADD_5.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6]|qx_net  ),
	. ci ( \carry_9_9__ADD_5|co_net  ),
	. co ( \carry_9_9__ADD_6|co_net  ),
	. s ( \carry_9_9__ADD_6|s_net  )
);
defparam carry_9_9__ADD_6.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_6.a_inv = "true";
defparam carry_9_9__ADD_6.PCK_LOCATION = "C18R13.lp0.add2.add0";
LUT6 ii3341 (
	. xy ( \ii3341|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii3341.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.lut_0";
defparam ii3341.PCK_LOCATION = "C6R14.lp0.lut_0";
defparam ii3341.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
SIO io_rx_decode_hsync_inst (
	. f_id ( )
,
	. clk_en ( ),
	. fclk ( ),
	. od ( {
		/* od [1] (nc) */ nc459 ,
		/* od [0] */ \ii2113|xy_net 
	} ),
	. oen ( ),
	. rstn ( ),
	. setn ( ),
	. PAD ( rx_decode_hsync )
);
defparam io_rx_decode_hsync_inst.DDR_PREG_EN = 0;
defparam io_rx_decode_hsync_inst.FCLK_GATE_EN = 0;
defparam io_rx_decode_hsync_inst.FOEN_SEL = 0;
defparam io_rx_decode_hsync_inst.RSTN_SYNC = 0;
defparam io_rx_decode_hsync_inst.OUT_SEL = 2;
defparam io_rx_decode_hsync_inst.DDR_EN = 0;
defparam io_rx_decode_hsync_inst.NDR = 15;
defparam io_rx_decode_hsync_inst.VPCI_EN = 0;
defparam io_rx_decode_hsync_inst.ID_RSTN_EN = 0;
defparam io_rx_decode_hsync_inst.KEEP = 0;
defparam io_rx_decode_hsync_inst.PDR = 15;
defparam io_rx_decode_hsync_inst.SETN_INV = 0;
defparam io_rx_decode_hsync_inst.SETN_SYNC = 0;
defparam io_rx_decode_hsync_inst.FIN_SEL = 0;
defparam io_rx_decode_hsync_inst.ID_SETN_EN = 0;
defparam io_rx_decode_hsync_inst.DDR_REG_EN = 0;
defparam io_rx_decode_hsync_inst.FOUT_SEL = 0;
defparam io_rx_decode_hsync_inst.OEN_RSTN_EN = 0;
defparam io_rx_decode_hsync_inst.NS_LV = 3;
defparam io_rx_decode_hsync_inst.optional_function = "";
defparam io_rx_decode_hsync_inst.OD_RSTN_EN = 0;
defparam io_rx_decode_hsync_inst.RSTN_INV = 0;
defparam io_rx_decode_hsync_inst.is_clk_io = "false";
defparam io_rx_decode_hsync_inst.PLACE_LOCATION = "C24R17.io_guts.iob_ck.I0.I60.Iioc0";
defparam io_rx_decode_hsync_inst.OEN_SETN_EN = 0;
defparam io_rx_decode_hsync_inst.OEN_SEL = 1;
defparam io_rx_decode_hsync_inst.PCK_LOCATION = "NONE";
defparam io_rx_decode_hsync_inst.OD_SETN_EN = 0;
defparam io_rx_decode_hsync_inst.CLK_INV = 0;
defparam io_rx_decode_hsync_inst.is_signal_monitor_io = 1'b0;
defparam io_rx_decode_hsync_inst.DDR_NREG_EN = 0;
defparam io_rx_decode_hsync_inst.RX_DIG_EN = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17]|qx_net  ),
	. di ( \ii2162|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17] .always_en = 0;
ADD1_A carry_12_0__ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6]|qx_net  ),
	. ci ( \carry_12_0__ADD_5|co_net  ),
	. co ( \carry_12_0__ADD_6|co_net  ),
	. s ( \carry_12_0__ADD_6|s_net  )
);
defparam carry_12_0__ADD_6.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_6.a_inv = "false";
defparam carry_12_0__ADD_6.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7]|qx_net  ),
	. ci ( \carry_9_9__ADD_6|co_net  ),
	. co ( \carry_9_9__ADD_7|co_net  ),
	. s ( \carry_9_9__ADD_7|s_net  )
);
defparam carry_9_9__ADD_7.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_7.a_inv = "true";
defparam carry_9_9__ADD_7.PCK_LOCATION = "C18R13.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .PCK_LOCATION = "C14R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[1] .always_en = 1;
LUT6 ii3342 (
	. xy ( \ii3342|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[8]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[0]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[8]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[0]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3342.PLACE_LOCATION = "C4R12.le_tile.le_guts.lp0.lut_0";
defparam ii3342.PCK_LOCATION = "C4R12.lp0.lut_0";
defparam ii3342.config_data = 64'b1111111110101010010101010000000011100100111001001110010011100100;
ADD1_A carry_12_0__ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7]|qx_net  ),
	. ci ( \carry_12_0__ADD_6|co_net  ),
	. co ( \carry_12_0__ADD_7|co_net  ),
	. s ( \carry_12_0__ADD_7|s_net  )
);
defparam carry_12_0__ADD_7.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_7.a_inv = "false";
defparam carry_12_0__ADD_7.PCK_LOCATION = "C8R4.lp0.add2.add0";
ADD1_A carry_9_9__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_9__ADD_7|co_net  ),
	. co ( \carry_9_9__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_9__ADD_8.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_9__ADD_8.a_inv = "false";
defparam carry_9_9__ADD_8.PCK_LOCATION = "C18R14.lp0.add2.add0";
LUT6 ii3343 (
	. xy ( \ii3343|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[24]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[16]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[24]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[16]_net  )
);
defparam ii3343.PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.lut_0";
defparam ii3343.PCK_LOCATION = "C4R13.lp0.lut_0";
defparam ii3343.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[14]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[14]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[14] .always_en = 1;
ADD1_A carry_12_0__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8]|qx_net  ),
	. ci ( \carry_12_0__ADD_7|co_net  ),
	. co ( \carry_12_0__ADD_8|co_net  ),
	. s ( \carry_12_0__ADD_8|s_net  )
);
defparam carry_12_0__ADD_8.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_8.a_inv = "false";
defparam carry_12_0__ADD_8.PCK_LOCATION = "C8R5.lp0.add2.add0";
LUT6 ii3344 (
	. xy ( \ii3344|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3343|xy_net  ),
	. f0 ( \ii3342|xy_net  )
);
defparam ii3344.PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.lut_0";
defparam ii3344.PCK_LOCATION = "C4R15.lp0.lut_0";
defparam ii3344.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
ADD1_A carry_12_0__ADD_9 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9]|qx_net  ),
	. ci ( \carry_12_0__ADD_8|co_net  ),
	. co ( \carry_12_0__ADD_9|co_net  ),
	. s ( \carry_12_0__ADD_9|s_net  )
);
defparam carry_12_0__ADD_9.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_9.a_inv = "false";
defparam carry_12_0__ADD_9.PCK_LOCATION = "C8R5.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0] .always_en = 1;
LUT6 ii3345 (
	. xy ( \ii3345|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[9]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[1]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[9]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[1]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3345.PLACE_LOCATION = "C4R12.le_tile.le_guts.lp0.lut_0";
defparam ii3345.PCK_LOCATION = "C4R12.lp0.lut_0";
defparam ii3345.config_data = 64'b1111111110101010010101010000000011100100111001001110010011100100;
REG \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3]|qx_net  ),
	. di ( \ii3386|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3] .always_en = 0;
LUT6 ii3346 (
	. xy ( \ii3346|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[25]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[17]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[25]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[17]_net  )
);
defparam ii3346.PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.lut_0";
defparam ii3346.PCK_LOCATION = "C4R13.lp0.lut_0";
defparam ii3346.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[8]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .PLACE_LOCATION = "C18R29.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .PCK_LOCATION = "C18R29.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3] .always_en = 1;
LUT6 ii3347 (
	. xy ( \ii3347|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3346|xy_net  ),
	. f0 ( \ii3345|xy_net  )
);
defparam ii3347.PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.lut_0";
defparam ii3347.PCK_LOCATION = "C4R15.lp0.lut_0";
defparam ii3347.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3] .always_en = 1;
LUT6 ii3348 (
	. xy ( \ii3348|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[2]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[10]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[2]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[10]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3348.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam ii3348.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam ii3348.config_data = 64'b1111111101010101101010100000000011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3]|qx_net  ),
	. di ( \ii2372|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .PCK_LOCATION = "C16R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2]|qx_net  ),
	. di ( \ii2243|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2] .always_en = 0;
LUT6 ii3349 (
	. xy ( \ii3349|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[26]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[18]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[26]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[18]_net  )
);
defparam ii3349.PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.lut_0";
defparam ii3349.PCK_LOCATION = "C4R13.lp0.lut_0";
defparam ii3349.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
LUT6 ii3350 (
	. xy ( \ii3350|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3349|xy_net  ),
	. f0 ( \ii3348|xy_net  )
);
defparam ii3350.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii3350.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii3350.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
REG \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1]|qx_net  ),
	. di ( \ii3368|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .PCK_LOCATION = "C4R16.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4]|qx_net  ),
	. di ( \ii2572|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1]|qx_net  ),
	. di ( \ii2432|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1] .always_en = 1;
REG \glue_cmd_s_reg[7]  (
	. qx ( \glue_cmd_s_reg[7]|qx_net  ),
	. di ( \mcu_arbiter_u_pfifo_u_inst|dout[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_cmd_s_reg[7] .latch_mode = 0;
defparam \glue_cmd_s_reg[7] .init = 0;
defparam \glue_cmd_s_reg[7] .PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.reg0";
defparam \glue_cmd_s_reg[7] .sr_inv = 1;
defparam \glue_cmd_s_reg[7] .sync_mode = 0;
defparam \glue_cmd_s_reg[7] .no_sr = 0;
defparam \glue_cmd_s_reg[7] .sr_value = 0;
defparam \glue_cmd_s_reg[7] .PCK_LOCATION = "C14R29.lp0.reg0";
defparam \glue_cmd_s_reg[7] .clk_inv = 0;
defparam \glue_cmd_s_reg[7] .en_inv = 0;
defparam \glue_cmd_s_reg[7] .always_en = 0;
LUT6 ii3351 (
	. xy ( \ii3351|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[3]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[11]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[3]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[11]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3351.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3351.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3351.config_data = 64'b1111111101010101101010100000000011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18]|qx_net  ),
	. di ( \ii2163|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .PCK_LOCATION = "C14R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[2] .always_en = 1;
LUT6 ii3352 (
	. xy ( \ii3352|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[27]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[19]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[27]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[19]_net  )
);
defparam ii3352.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3352.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3352.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
LUT6 ii3353 (
	. xy ( \ii3353|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3352|xy_net  ),
	. f0 ( \ii3351|xy_net  )
);
defparam ii3353.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii3353.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii3353.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[15]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[15]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[15] .always_en = 1;
LUT6 ii3354 (
	. xy ( \ii3354|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[4]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[12]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[4]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[12]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3354.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3354.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3354.config_data = 64'b1111111101010101101010100000000011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .PLACE_LOCATION = "C8R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .PCK_LOCATION = "C8R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1] .always_en = 1;
LUT6 ii3355 (
	. xy ( \ii3355|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[28]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[20]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[28]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[20]_net  )
);
defparam ii3355.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3355.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3355.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
REG \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4]|qx_net  ),
	. di ( \ii3386|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4] .always_en = 0;
LUT6 ii3356 (
	. xy ( \ii3356|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3355|xy_net  ),
	. f0 ( \ii3354|xy_net  )
);
defparam ii3356.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii3356.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii3356.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2000 (
	. xy ( \ii2000|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8]|qx_net  )
);
defparam ii2000.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.lut_0";
defparam ii2000.PCK_LOCATION = "C20R23.lp0.lut_0";
defparam ii2000.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii3357 (
	. xy ( \ii3357|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[5]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[13]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[5]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[13]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3357.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3357.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3357.config_data = 64'b1111111101010101101010100000000011011000110110001101100011011000;
REG uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg (
	. qx ( \uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd_valid_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.latch_mode = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.init = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.sr_inv = 1;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.sync_mode = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.no_sr = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.sr_value = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.PCK_LOCATION = "C4R7.lp0.reg0";
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.clk_inv = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.en_inv = 0;
defparam uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4] .always_en = 1;
LUT6 ii2001 (
	. xy ( \ii2001|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9]|qx_net  )
);
defparam ii2001.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.lut_0";
defparam ii2001.PCK_LOCATION = "C20R23.lp0.lut_0";
defparam ii2001.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii3358 (
	. xy ( \ii3358|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[29]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[21]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[29]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[21]_net  )
);
defparam ii3358.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3358.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3358.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4]|qx_net  ),
	. di ( \ii2373|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3]|qx_net  ),
	. di ( \ii2246|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3] .always_en = 0;
LUT6 ii3359 (
	. xy ( \ii3359|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3358|xy_net  ),
	. f0 ( \ii3357|xy_net  )
);
defparam ii3359.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii3359.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii3359.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii3360 (
	. xy ( \ii3360|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[6]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[14]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[6]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[14]_net  )
);
defparam ii3360.PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.lut_0";
defparam ii3360.PCK_LOCATION = "C4R13.lp0.lut_0";
defparam ii3360.config_data = 64'b1111111100000000110011001100110011110000111100001010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5]|qx_net  ),
	. di ( \ii2573|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2]|qx_net  ),
	. di ( \ii2433|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2] .always_en = 1;
LUT6 ii3361 (
	. xy ( \ii3361|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[30]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[22]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[30]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[22]_net  )
);
defparam ii3361.PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.lut_0";
defparam ii3361.PCK_LOCATION = "C4R13.lp0.lut_0";
defparam ii3361.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20]|qx_net  ),
	. di ( \ii2168|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19]|qx_net  ),
	. di ( \ii2164|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .PCK_LOCATION = "C14R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[3] .always_en = 1;
LUT6 ii3362 (
	. xy ( \ii3362|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3361|xy_net  ),
	. f0 ( \ii3360|xy_net  )
);
defparam ii3362.PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.lut_0";
defparam ii3362.PCK_LOCATION = "C4R15.lp0.lut_0";
defparam ii3362.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
REG glue_rx_packet_tx_packet_rx_hsync_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. di ( \ii2294|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_hsync_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_hsync_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.PCK_LOCATION = "C10R5.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_hsync_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_hsync_reg.always_en = 1;
LUT6 ii3363 (
	. xy ( \ii3363|xy_net  ),
	. f5 ( \mipi_inst_u_mipi2|pready_net  ),
	. f4 ( \mipi_inst_u_mipi2|prdata[7]_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[15]_net  ),
	. f2 ( \mipi_inst_u_mipi1|prdata[7]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[15]_net  ),
	. f0 ( \ii3341|xy_net  )
);
defparam ii3363.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3363.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3363.config_data = 64'b1111111101010101101010100000000011011000110110001101100011011000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[16]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[16]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[16] .always_en = 1;
LUT6 ii3364 (
	. xy ( \ii3364|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f4 ( \mipi_inst_u_mipi2|pready_net  ),
	. f3 ( \mipi_inst_u_mipi2|prdata[31]_net  ),
	. f2 ( \mipi_inst_u_mipi2|prdata[23]_net  ),
	. f1 ( \mipi_inst_u_mipi1|prdata[31]_net  ),
	. f0 ( \mipi_inst_u_mipi1|prdata[23]_net  )
);
defparam ii3364.PLACE_LOCATION = "C6R13.le_tile.le_guts.lp0.lut_0";
defparam ii3364.PCK_LOCATION = "C6R13.lp0.lut_0";
defparam ii3364.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2] .always_en = 1;
LUT6 ii3365 (
	. xy ( \ii3365|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \ii3364|xy_net  ),
	. f0 ( \ii3363|xy_net  )
);
defparam ii3365.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii3365.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii3365.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
REG \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5]|qx_net  ),
	. di ( \ii3387|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3381|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .PCK_LOCATION = "C6R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5] .always_en = 0;
LUT6 ii3366 (
	. xy ( \ii3366|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memwr_comb_net  ),
	. f0 ( \ii3317|xy_net  )
);
defparam ii3366.PLACE_LOCATION = "C8R17.le_tile.le_guts.lp0.lut_0";
defparam ii3366.PCK_LOCATION = "C8R17.lp0.lut_0";
defparam ii3366.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii3367 (
	. xy ( \ii3367|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0]|qx_net  )
);
defparam ii3367.PLACE_LOCATION = "C4R17.le_tile.le_guts.lp0.lut_0";
defparam ii3367.PCK_LOCATION = "C4R17.lp0.lut_0";
defparam ii3367.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5] .always_en = 1;
LUT6 ii3368 (
	. xy ( \ii3368|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[1]|qx_net  ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_byte_cnt_reg[0]|qx_net  )
);
defparam ii3368.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.lut_0";
defparam ii3368.PCK_LOCATION = "C4R16.lp0.lut_0";
defparam ii3368.config_data = 64'b0110011001100110011001100110011001100110011001100110011001100110;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5]|qx_net  ),
	. di ( \ii2374|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4]|qx_net  ),
	. di ( \ii2247|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4] .always_en = 0;
REG glue_rx_packet_tx_packet_u_scaler_t47_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.PLACE_LOCATION = "C20R24.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.PCK_LOCATION = "C20R24.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t47_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_5__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[0] .always_en = 1;
LUT6 ii3369 (
	. xy ( \ii3369|xy_net  ),
	. f5 ( ),
	. f4 ( \u_8051_u_h6_8051|memrd_comb_net  ),
	. f3 ( \u_8051_u_h6_8051|mempsrd_comb_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[17]_net  ),
	. f1 ( \ii2047|xy_net  ),
	. f0 ( \ii2046|xy_net  )
);
defparam ii3369.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.lut_0";
defparam ii3369.PCK_LOCATION = "C4R18.lp0.lut_0";
defparam ii3369.config_data = 64'b0101010100010101010101010001000101010101000101010101010100010001;
LUT6 ii3370 (
	. xy ( \ii3370|xy_net  ),
	. f5 ( ),
	. f4 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15]|qx_net  ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12]|qx_net  ),
	. f0 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11]|qx_net  )
);
defparam ii3370.PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.lut_0";
defparam ii3370.PCK_LOCATION = "C4R6.lp0.lut_0";
defparam ii3370.config_data = 64'b0000100000000000000000000000000000001000000000000000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6]|qx_net  ),
	. di ( \ii2574|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .PCK_LOCATION = "C18R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3]|qx_net  ),
	. di ( \ii2434|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .PCK_LOCATION = "C10R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3] .always_en = 1;
LUT6 ii3371 (
	. xy ( \ii3371|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  ),
	. f0 ( \ii3370|xy_net  )
);
defparam ii3371.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3371.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3371.config_data = 64'b0000001000000000000000100000000000000010000000000000001000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21]|qx_net  ),
	. di ( \ii2169|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .PCK_LOCATION = "C14R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[4] .always_en = 1;
LUT6 ii3372 (
	. xy ( \ii3372|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13]|qx_net  ),
	. f0 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12]|qx_net  )
);
defparam ii3372.PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.lut_0";
defparam ii3372.PCK_LOCATION = "C4R6.lp0.lut_0";
defparam ii3372.config_data = 64'b0010000000000000001000000000000000100000000000000010000000000000;
LUT6 ii3373 (
	. xy ( \ii3373|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[11]|qx_net  ),
	. f0 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  )
);
defparam ii3373.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3373.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3373.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[17]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[17]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[17] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t16_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.PCK_LOCATION = "C18R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t16_out1_reg.always_en = 1;
LUT6 ii3374 (
	. xy ( \ii3374|xy_net  ),
	. f5 ( ),
	. f4 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f2 ( \ii3373|xy_net  ),
	. f1 ( \ii3372|xy_net  ),
	. f0 ( \ii3371|xy_net  )
);
defparam ii3374.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3374.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3374.config_data = 64'b0101010101010101010101010001010101010101010101010101010100010101;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0]|qx_net  ),
	. di ( \ii2511|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .PLACE_LOCATION = "C8R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .PCK_LOCATION = "C8R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3] .always_en = 1;
LUT6 ii3375 (
	. xy ( \ii3375|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  ),
	. f0 ( \ii3370|xy_net  )
);
defparam ii3375.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3375.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3375.config_data = 64'b0010000000100000001000000010000000100000001000000010000000100000;
LUT6 ii3376 (
	. xy ( \ii3376|xy_net  ),
	. f5 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[5]|qx_net  ),
	. f4 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[4]|qx_net  ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[3]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[2]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[1]|qx_net  ),
	. f0 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[0]|qx_net  )
);
defparam ii3376.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii3376.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii3376.config_data = 64'b0000000000000000000000000000000000000000000100000000000001000000;
LUT6 ii3377 (
	. xy ( \ii3377|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_valid_d_reg|qx_net  ),
	. f0 ( \ii3376|xy_net  )
);
defparam ii3377.PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.lut_0";
defparam ii3377.PCK_LOCATION = "C6R6.lp0.lut_0";
defparam ii3377.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[22]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf.PLACE_LOCATION = "C8R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf.PCK_LOCATION = "C8R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6] .always_en = 1;
LUT6 ii3378 (
	. xy ( \ii3378|xy_net  ),
	. f5 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f4 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[15]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[14]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[13]|qx_net  ),
	. f0 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[12]|qx_net  )
);
defparam ii3378.PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.lut_0";
defparam ii3378.PCK_LOCATION = "C4R6.lp0.lut_0";
defparam ii3378.config_data = 64'b0000100000000000000000000000000000000000000000000000000000000000;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6]|qx_net  ),
	. di ( \ii2375|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5]|qx_net  ),
	. di ( \ii2248|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5] .always_en = 0;
ADD1_A carry_9_11__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_11__ADD_0|co_net  ),
	. s ( \carry_9_11__ADD_0|s_net  )
);
defparam carry_9_11__ADD_0.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_0.a_inv = "true";
defparam carry_9_11__ADD_0.PCK_LOCATION = "C20R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_5__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[1] .always_en = 1;
LUT6 ii3379 (
	. xy ( \ii3379|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f0 ( \ii3378|xy_net  )
);
defparam ii3379.PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.lut_0";
defparam ii3379.PCK_LOCATION = "C6R6.lp0.lut_0";
defparam ii3379.config_data = 64'b0101010001010100010101000101010001010100010101000101010001010100;
LUT6 ii3380 (
	. xy ( \ii3380|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f0 ( \ii3372|xy_net  )
);
defparam ii3380.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3380.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3380.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7]|qx_net  ),
	. di ( \ii2575|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4]|qx_net  ),
	. di ( \ii2435|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4] .always_en = 1;
ADD1_A carry_9_11__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1]|qx_net  ),
	. ci ( \carry_9_11__ADD_0|co_net  ),
	. co ( \carry_9_11__ADD_1|co_net  ),
	. s ( \carry_9_11__ADD_1|s_net  )
);
defparam carry_9_11__ADD_1.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_1.a_inv = "true";
defparam carry_9_11__ADD_1.PCK_LOCATION = "C20R8.lp0.add2.add0";
LUT6 ii3381 (
	. xy ( \ii3381|xy_net  ),
	. f5 ( ),
	. f4 ( \ii3373|xy_net  ),
	. f3 ( \ii3380|xy_net  ),
	. f2 ( \ii3379|xy_net  ),
	. f1 ( \ii3377|xy_net  ),
	. f0 ( \ii3375|xy_net  )
);
defparam ii3381.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3381.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3381.config_data = 64'b1000100010001100100010001000100010001000100011001000100010001000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22]|qx_net  ),
	. di ( \ii2170|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22] .always_en = 0;
ADD1_A carry_9_11__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2]|qx_net  ),
	. ci ( \carry_9_11__ADD_1|co_net  ),
	. co ( \carry_9_11__ADD_2|co_net  ),
	. s ( \carry_9_11__ADD_2|s_net  )
);
defparam carry_9_11__ADD_2.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_2.a_inv = "true";
defparam carry_9_11__ADD_2.PCK_LOCATION = "C20R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .PCK_LOCATION = "C10R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_In1p_reg[5] .always_en = 1;
LUT6 ii3382 (
	. xy ( \ii3382|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  ),
	. f0 ( \ii3370|xy_net  )
);
defparam ii3382.PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.lut_0";
defparam ii3382.PCK_LOCATION = "C6R6.lp0.lut_0";
defparam ii3382.config_data = 64'b0010000000001000001000000000100000100000000010000010000000001000;
ADD1_A carry_9_11__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3]|qx_net  ),
	. ci ( \carry_9_11__ADD_2|co_net  ),
	. co ( \carry_9_11__ADD_3|co_net  ),
	. s ( \carry_9_11__ADD_3|s_net  )
);
defparam carry_9_11__ADD_3.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_3.a_inv = "true";
defparam carry_9_11__ADD_3.PCK_LOCATION = "C20R8.lp0.add2.add0";
LUT6 ii3383 (
	. xy ( \ii3383|xy_net  ),
	. f5 ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1]|qx_net  ),
	. f4 ( \ii3378|xy_net  ),
	. f3 ( \ii3373|xy_net  ),
	. f2 ( \ii3382|xy_net  ),
	. f1 ( \ii3377|xy_net  ),
	. f0 ( \ii3371|xy_net  )
);
defparam ii3383.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3383.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3383.config_data = 64'b1011111110111111101111111011111110001100100010001000100010001000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[18]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[18]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[18] .always_en = 1;
ADD1_A carry_9_11__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4]|qx_net  ),
	. ci ( \carry_9_11__ADD_3|co_net  ),
	. co ( \carry_9_11__ADD_4|co_net  ),
	. s ( \carry_9_11__ADD_4|s_net  )
);
defparam carry_9_11__ADD_4.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_4.a_inv = "true";
defparam carry_9_11__ADD_4.PCK_LOCATION = "C20R8.lp0.add2.add0";
LUT6 ii2026 (
	. xy ( \ii2026|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2026.PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.lut_0";
defparam ii2026.PCK_LOCATION = "C18R16.lp0.lut_0";
defparam ii2026.config_data = 64'b1000000011000000100010001100110010000000110000001000100011001100;
LUT6 ii3384 (
	. xy ( \ii3384|xy_net  ),
	. f5 ( \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4]|qx_net  ),
	. f4 ( \ii3373|xy_net  ),
	. f3 ( \ii3380|xy_net  ),
	. f2 ( \ii3379|xy_net  ),
	. f1 ( \ii3377|xy_net  ),
	. f0 ( \ii3375|xy_net  )
);
defparam ii3384.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3384.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3384.config_data = 64'b1111111111111011111111111111111110001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1]|qx_net  ),
	. di ( \ii2512|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1] .always_en = 1;
ADD1_A carry_9_11__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5]|qx_net  ),
	. ci ( \carry_9_11__ADD_4|co_net  ),
	. co ( \carry_9_11__ADD_5|co_net  ),
	. s ( \carry_9_11__ADD_5|s_net  )
);
defparam carry_9_11__ADD_5.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_5.a_inv = "true";
defparam carry_9_11__ADD_5.PCK_LOCATION = "C20R8.lp0.add2.add0";
LUT6 ii2027 (
	. xy ( \ii2027|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_1|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2027.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2027.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2027.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
LUT6 ii3385 (
	. xy ( \ii3385|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f0 ( \ii3375|xy_net  )
);
defparam ii3385.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3385.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3385.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
ADD1_A carry_9_11__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6]|qx_net  ),
	. ci ( \carry_9_11__ADD_5|co_net  ),
	. co ( \carry_9_11__ADD_6|co_net  ),
	. s ( \carry_9_11__ADD_6|s_net  )
);
defparam carry_9_11__ADD_6.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_6.a_inv = "true";
defparam carry_9_11__ADD_6.PCK_LOCATION = "C20R8.lp0.add2.add0";
LUT6 ii2028 (
	. xy ( \ii2028|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_2|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2028.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2028.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2028.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
LUT6 ii3386 (
	. xy ( \ii3386|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[9]|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[8]|qx_net  ),
	. f1 ( \uut_dataReadBack_mipi_periph_rx_cmd_d_reg[10]|qx_net  ),
	. f0 ( \ii3370|xy_net  )
);
defparam ii3386.PLACE_LOCATION = "C6R5.le_tile.le_guts.lp0.lut_0";
defparam ii3386.PCK_LOCATION = "C6R5.lp0.lut_0";
defparam ii3386.config_data = 64'b1101110111110111110111011111011111011101111101111101110111110111;
ADD1_A carry_9_11__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7]|qx_net  ),
	. ci ( \carry_9_11__ADD_6|co_net  ),
	. co ( \carry_9_11__ADD_7|co_net  ),
	. s ( \carry_9_11__ADD_7|s_net  )
);
defparam carry_9_11__ADD_7.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_7.a_inv = "true";
defparam carry_9_11__ADD_7.PCK_LOCATION = "C20R8.lp0.add2.add0";
LUT6 ii2029 (
	. xy ( \ii2029|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_3|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2029.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2029.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2029.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
LUT6 ii2030 (
	. xy ( \ii2030|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_4|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2030.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2030.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2030.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
LUT6 ii3387 (
	. xy ( \ii3387|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \ii3386|xy_net  )
);
defparam ii3387.PLACE_LOCATION = "C6R4.le_tile.le_guts.lp0.lut_0";
defparam ii3387.PCK_LOCATION = "C6R4.lp0.lut_0";
defparam ii3387.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
REG \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d0|doa[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7] .always_en = 1;
ADD1_A carry_9_11__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_11__ADD_7|co_net  ),
	. co ( \carry_9_11__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_11__ADD_8.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_11__ADD_8.a_inv = "false";
defparam carry_9_11__ADD_8.PCK_LOCATION = "C20R9.lp0.add2.add0";
LUT6 ii2031 (
	. xy ( \ii2031|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_5|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2031.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2031.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2031.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
LUT6 ii3388 (
	. xy ( \ii3388|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \uut_dataReadBack_mipi_periph_tx_cmd_req_reg|qx_net  ),
	. f2 ( \uut_dataReadBack_mipi_periph_dphy_direction_d_reg|qx_net  ),
	. f1 ( \mipi_inst_u_mipi1|periph_tx_cmd_ack_net  ),
	. f0 ( \mipi_inst_u_mipi1|periph_dphy_direction_net  )
);
defparam ii3388.PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.lut_0";
defparam ii3388.PCK_LOCATION = "C4R7.lp0.lut_0";
defparam ii3388.config_data = 64'b0111001101010000011100110101000001110011010100000111001101010000;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7]|qx_net  ),
	. di ( \ii2376|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6]|qx_net  ),
	. di ( \ii2249|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_5__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[2] .always_en = 1;
LUT6 ii2032 (
	. xy ( \ii2032|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_6|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2032.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2032.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2032.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8]|qx_net  ),
	. di ( \ii2576|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5]|qx_net  ),
	. di ( \ii2436|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5] .always_en = 1;
LUT6 ii2033 (
	. xy ( \ii2033|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \carry_11_ADD_7|s_net  ),
	. f1 ( \ii1982_dup|xy_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2033.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.lut_0";
defparam ii2033.PCK_LOCATION = "C20R16.lp0.lut_0";
defparam ii2033.config_data = 64'b1100100000000000110010001100100011001000000000001100100011001000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23]|qx_net  ),
	. di ( \ii2171|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23] .always_en = 0;
LUT6 ii2034 (
	. xy ( \ii2034|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \ii1982_dup|xy_net  ),
	. f1 ( \carry_11_ADD_8|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2034.PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.lut_0";
defparam ii2034.PCK_LOCATION = "C18R16.lp0.lut_0";
defparam ii2034.config_data = 64'b1110000000000000111000001110000011100000000000001110000011100000;
LUT6 ii2035 (
	. xy ( \ii2035|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f2 ( \ii1982_dup|xy_net  ),
	. f1 ( \carry_11_ADD_9|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2035.PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.lut_0";
defparam ii2035.PCK_LOCATION = "C18R16.lp0.lut_0";
defparam ii2035.config_data = 64'b1110000000000000111000001110000011100000000000001110000011100000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[19]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[19]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[19] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[20]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[20]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[20] .always_en = 1;
LUT6 ii2036 (
	. xy ( \ii2036|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rd_cmd_flag_reg|qx_net  ),
	. f0 ( \mipi_inst_u_mipi2|host_tx_payload_en_net  )
);
defparam ii2036.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2036.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2036.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2]|qx_net  ),
	. di ( \ii2513|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[10] .always_en = 1;
LUT6 ii2037 (
	. xy ( \ii2037|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \mcu_arbiter_fifo_clr_s_reg|qx_net  ),
	. f1 ( \mcu_arbiter_fifo_clr_d_reg|qx_net  ),
	. f0 ( \ii1982_dup|xy_net  )
);
defparam ii2037.PLACE_LOCATION = "C4R24.le_tile.le_guts.lp0.lut_0";
defparam ii2037.PCK_LOCATION = "C4R24.lp0.lut_0";
defparam ii2037.config_data = 64'b1000101010001010100010101000101010001010100010101000101010001010;
LUT6 ii2038 (
	. xy ( \ii2038|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[17]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[11]_net  )
);
defparam ii2038.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.lut_0";
defparam ii2038.PCK_LOCATION = "C4R18.lp0.lut_0";
defparam ii2038.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii2039 (
	. xy ( \ii2039|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \u_8051_u_h6_8051|memwr_comb_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[3]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \ii2038|xy_net  )
);
defparam ii2039.PLACE_LOCATION = "C4R17.le_tile.le_guts.lp0.lut_0";
defparam ii2039.PCK_LOCATION = "C4R17.lp0.lut_0";
defparam ii2039.config_data = 64'b0000001000000000000000100000000000000010000000000000001000000000;
LUT6 ii2040 (
	. xy ( \ii2040|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \mcu_arbiter_fifo_wr_d_reg|qx_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[2]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f0 ( \ii2039|xy_net  )
);
defparam ii2040.PLACE_LOCATION = "C4R19.le_tile.le_guts.lp0.lut_0";
defparam ii2040.PCK_LOCATION = "C4R19.lp0.lut_0";
defparam ii2040.config_data = 64'b1111111111111101111111111111110111111111111111011111111111111101;
LUT6 ii2041 (
	. xy ( \ii2041|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  )
);
defparam ii2041.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2041.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2041.config_data = 64'b1110111011101110111011101110111011101110111011101110111011101110;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8]|qx_net  ),
	. di ( \ii2377|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7]|qx_net  ),
	. di ( \ii2250|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_5__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[3] .always_en = 1;
LUT6 ii2042 (
	. xy ( \ii2042|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f0 ( \ii2041|xy_net  )
);
defparam ii2042.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2042.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2042.config_data = 64'b1101111111011111110111111101111111011111110111111101111111011111;
REG \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9]|qx_net  ),
	. di ( \ii2577|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6]|qx_net  ),
	. di ( \ii2437|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6] .always_en = 1;
LUT6 ii2043 (
	. xy ( \ii2043|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f0 ( \ii2041|xy_net  )
);
defparam ii2043.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2043.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2043.config_data = 64'b1101111111011111110111111101111111011111110111111101111111011111;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24]|qx_net  ),
	. di ( \ii2172|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24] .always_en = 0;
LUT6 ii2044 (
	. xy ( \ii2044|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. f0 ( \ii2041|xy_net  )
);
defparam ii2044.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.lut_0";
defparam ii2044.PCK_LOCATION = "C6R20.lp0.lut_0";
defparam ii2044.config_data = 64'b0111110101111101011111010111110101111101011111010111110101111101;
LUT6 ii2045 (
	. xy ( \ii2045|xy_net  ),
	. f5 ( \u_8051_u_h6_8051|memaddr_comb[20]_net  ),
	. f4 ( \u_8051_u_h6_8051|memaddr_comb[22]_net  ),
	. f3 ( \u_8051_u_h6_8051|memaddr_comb[15]_net  ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[17]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[19]_net  ),
	. f0 ( \u_8051_u_h6_8051|memaddr_comb[21]_net  )
);
defparam ii2045.PLACE_LOCATION = "C6R16.le_tile.le_guts.lp0.lut_0";
defparam ii2045.PCK_LOCATION = "C6R16.lp0.lut_0";
defparam ii2045.config_data = 64'b0000000000000000000000000000000000000000000000000000000000000001;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[12]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf.PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf.PCK_LOCATION = "C14R13.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[21]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[21]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[21] .always_en = 1;
LUT6 ii2046 (
	. xy ( \ii2046|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[16]_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[18]_net  ),
	. f0 ( \ii2045|xy_net  )
);
defparam ii2046.PLACE_LOCATION = "C6R19.le_tile.le_guts.lp0.lut_0";
defparam ii2046.PCK_LOCATION = "C6R19.lp0.lut_0";
defparam ii2046.config_data = 64'b1111110111111101111111011111110111111101111111011111110111111101;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3]|qx_net  ),
	. di ( \ii2514|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[11] .always_en = 1;
LUT6 ii2047 (
	. xy ( \ii2047|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \u_8051_u_h6_8051|memaddr_comb[17]_net  ),
	. f1 ( \u_8051_u_h6_8051|memwr_comb_net  ),
	. f0 ( \u_8051_u_h6_8051|mempswr_comb_net  )
);
defparam ii2047.PLACE_LOCATION = "C4R19.le_tile.le_guts.lp0.lut_0";
defparam ii2047.PCK_LOCATION = "C4R19.lp0.lut_0";
defparam ii2047.config_data = 64'b0101000101010001010100010101000101010001010100010101000101010001;
REG glue_rx_packet_tx_packet_u_scaler_t75_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t75_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.PCK_LOCATION = "C8R20.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t75_out1_reg.always_en = 1;
LUT6 ii2048 (
	. xy ( \ii2048|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \mcu_arbiter_func_reg[0]|qx_net  ),
	. f1 ( \u_8051_u_h6_8051|port0o[2]_net  ),
	. f0 ( \ii1982_dup|xy_net  )
);
defparam ii2048.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam ii2048.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam ii2048.config_data = 64'b1000000010000000100000001000000010000000100000001000000010000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[0] .always_en = 1;
LUT6 ii2049 (
	. xy ( \ii2049|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \ii2048|xy_net  )
);
defparam ii2049.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii2049.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii2049.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 ii2050 (
	. xy ( \ii2050|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \mcu_arbiter_u_emif2apb_fpga_HRD_reg|qx_net  ),
	. f1 ( \u_8051_u_h6_8051|memaddr_comb[17]_net  ),
	. f0 ( \mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf|xy_net  )
);
defparam ii2050.PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.lut_0";
defparam ii2050.PCK_LOCATION = "C4R14.lp0.lut_0";
defparam ii2050.config_data = 64'b1100100011001000110010001100100011001000110010001100100011001000;
LUT6 ii2051 (
	. xy ( \ii2051|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_mipi_sel_reg|qx_net  ),
	. f0 ( \ii2050|xy_net  )
);
defparam ii2051.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2051.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2051.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9]|qx_net  ),
	. di ( \ii2378|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8]|qx_net  ),
	. di ( \ii2251|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_5__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[4] .always_en = 1;
LUT6 ii2052 (
	. xy ( \ii2052|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[0]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2052.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2052.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2052.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7]|qx_net  ),
	. di ( \ii2438|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7] .always_en = 1;
LUT6 ii2053 (
	. xy ( \ii2053|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[10]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2053.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2053.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2053.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25]|qx_net  ),
	. di ( \ii2173|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25] .always_en = 0;
LUT6 ii2054 (
	. xy ( \ii2054|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[11]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2054.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2054.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2054.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2055 (
	. xy ( \ii2055|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[12]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2055.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2055.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2055.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG mcu_arbiter_data_sel_reg (
	. qx ( \mcu_arbiter_data_sel_reg|qx_net  ),
	. di ( \ii3319|xy_net  ),
	. sr ( ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_data_sel_reg.latch_mode = 0;
defparam mcu_arbiter_data_sel_reg.init = 0;
defparam mcu_arbiter_data_sel_reg.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_data_sel_reg.sr_inv = 0;
defparam mcu_arbiter_data_sel_reg.sync_mode = 1;
defparam mcu_arbiter_data_sel_reg.no_sr = 1;
defparam mcu_arbiter_data_sel_reg.sr_value = 0;
defparam mcu_arbiter_data_sel_reg.PCK_LOCATION = "C4R18.lp0.reg0";
defparam mcu_arbiter_data_sel_reg.clk_inv = 0;
defparam mcu_arbiter_data_sel_reg.en_inv = 0;
defparam mcu_arbiter_data_sel_reg.always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[22]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[22]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[22] .always_en = 1;
LUT6 ii2056 (
	. xy ( \ii2056|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[13]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2056.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2056.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2056.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4]|qx_net  ),
	. di ( \ii2515|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t13_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.PCK_LOCATION = "C18R22.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t13_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[12] .always_en = 1;
LUT6 ii2057 (
	. xy ( \ii2057|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[14]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2057.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2057.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2057.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2058 (
	. xy ( \ii2058|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[15]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2058.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2058.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2058.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG glue_rx_packet_tx_packet_u_scaler_t105_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t105_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t71_out1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.PLACE_LOCATION = "C20R24.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.PCK_LOCATION = "C20R24.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t105_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[1] .always_en = 1;
LUT6 ii2059 (
	. xy ( \ii2059|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[1]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2059.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2059.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2059.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2060 (
	. xy ( \ii2060|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[2]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2060.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2060.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2060.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2061 (
	. xy ( \ii2061|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[3]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2061.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2061.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2061.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9]|qx_net  ),
	. di ( \ii2252|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_5__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[5] .always_en = 1;
LUT6 ii2062 (
	. xy ( \ii2062|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[4]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2062.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2062.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2062.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2063 (
	. xy ( \ii2063|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[5]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2063.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2063.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2063.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26]|qx_net  ),
	. di ( \ii2174|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26] .always_en = 0;
LUT6 ii2064 (
	. xy ( \ii2064|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[6]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2064.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2064.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2064.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG glue_rd_start_d_reg (
	. qx ( \glue_rd_start_d_reg|qx_net  ),
	. di ( \glue_rd_start_s_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rd_start_d_reg.latch_mode = 0;
defparam glue_rd_start_d_reg.init = 0;
defparam glue_rd_start_d_reg.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam glue_rd_start_d_reg.sr_inv = 1;
defparam glue_rd_start_d_reg.sync_mode = 0;
defparam glue_rd_start_d_reg.no_sr = 0;
defparam glue_rd_start_d_reg.sr_value = 0;
defparam glue_rd_start_d_reg.PCK_LOCATION = "C16R17.lp0.reg0";
defparam glue_rd_start_d_reg.clk_inv = 0;
defparam glue_rd_start_d_reg.en_inv = 0;
defparam glue_rd_start_d_reg.always_en = 1;
LUT6 ii2065 (
	. xy ( \ii2065|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[7]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2065.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2065.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2065.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[23]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[23]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[23] .always_en = 1;
LUT6 ii2066 (
	. xy ( \ii2066|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[8]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2066.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2066.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2066.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5]|qx_net  ),
	. di ( \ii2516|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[13] .always_en = 1;
LUT6 ii2067 (
	. xy ( \ii2067|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57]|qx_net  ),
	. f1 ( \glue_dnum_s_reg[9]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2067.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2067.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2067.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2068 (
	. xy ( \ii2068|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]|qx_net  ),
	. f1 ( \glue_cmd_s_reg[0]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2068.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.lut_0";
defparam ii2068.PCK_LOCATION = "C14R25.lp0.lut_0";
defparam ii2068.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[2] .always_en = 1;
LUT6 ii2069 (
	. xy ( \ii2069|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]|qx_net  ),
	. f1 ( \glue_cmd_s_reg[1]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2069.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2069.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2069.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2070 (
	. xy ( \ii2070|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]|qx_net  ),
	. f1 ( \glue_cmd_s_reg[2]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2070.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2070.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2070.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2071 (
	. xy ( \ii2071|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]|qx_net  ),
	. f1 ( \glue_cmd_s_reg[3]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2071.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2071.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2071.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_5__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[6] .always_en = 1;
LUT6 ii2072 (
	. xy ( \ii2072|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]|qx_net  ),
	. f1 ( \glue_cmd_s_reg[4]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2072.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2072.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2072.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG rstn_r_reg (
	. qx ( \rstn_r_reg|qx_net  ),
	. di ( \u_pll_pll_u0|PLOCK_net  ),
	. sr ( ),
	. en ( ),
	. clk ( \u_osc|OSC_net  )
);
defparam rstn_r_reg.latch_mode = 0;
defparam rstn_r_reg.init = 0;
defparam rstn_r_reg.PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam rstn_r_reg.sr_inv = 0;
defparam rstn_r_reg.sync_mode = 1;
defparam rstn_r_reg.no_sr = 1;
defparam rstn_r_reg.sr_value = 0;
defparam rstn_r_reg.PCK_LOCATION = "C20R17.lp0.reg0";
defparam rstn_r_reg.clk_inv = 0;
defparam rstn_r_reg.en_inv = 0;
defparam rstn_r_reg.always_en = 1;
LUT6 ii2073 (
	. xy ( \ii2073|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]|qx_net  ),
	. f1 ( \glue_cmd_s_reg[5]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2073.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2073.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2073.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27]|qx_net  ),
	. di ( \ii2175|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27] .always_en = 0;
LUT6 ii2074 (
	. xy ( \ii2074|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]|qx_net  )
);
defparam ii2074.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2074.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2074.config_data = 64'b0000000000000001000000000000000100000000000000010000000000000001;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10]|qx_net  ),
	. di ( \ii2557|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .PCK_LOCATION = "C20R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10] .always_en = 1;
LUT6 ii2075 (
	. xy ( \ii2075|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]|qx_net  ),
	. f0 ( \ii2074|xy_net  )
);
defparam ii2075.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2075.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2075.config_data = 64'b1111111111111111111111111111110111111111111111111111111111111101;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[24]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[24]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[24] .always_en = 1;
LUT6 ii2076 (
	. xy ( \ii2076|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg|qx_net  ),
	. f2 ( \glue_pasm_cmd_rq_o_reg|qx_net  ),
	. f1 ( \ii2075|xy_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2076.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2076.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2076.config_data = 64'b1101100001010000110110000101000011011000010100001101100001010000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6]|qx_net  ),
	. di ( \ii2517|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .PLACE_LOCATION = "C20R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .PCK_LOCATION = "C20R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[14] .always_en = 1;
LUT6 ii2077 (
	. xy ( \ii2077|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_cmd_s_reg[6]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2077.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.lut_0";
defparam ii2077.PCK_LOCATION = "C14R30.lp0.lut_0";
defparam ii2077.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10]|qx_net  ),
	. di ( \ii2368|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10] .always_en = 0;
LUT6 ii2078 (
	. xy ( \ii2078|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_cmd_s_reg[7]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2078.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.lut_0";
defparam ii2078.PCK_LOCATION = "C14R30.lp0.lut_0";
defparam ii2078.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .PCK_LOCATION = "C20R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[3] .always_en = 1;
LUT6 ii2079 (
	. xy ( \ii2079|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_func_reg[1]|qx_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2079.PLACE_LOCATION = "C10R23.le_tile.le_guts.lp0.lut_0";
defparam ii2079.PCK_LOCATION = "C10R23.lp0.lut_0";
defparam ii2079.config_data = 64'b1110111011101110111011101110111011101110111011101110111011101110;
LUT6 ii2080 (
	. xy ( \ii2080|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[0]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[0]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2080.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2080.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2080.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2081 (
	. xy ( \ii2081|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[10]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2081.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2081.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2081.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_5__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .PCK_LOCATION = "C14R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[7] .always_en = 1;
LUT6 ii1982 (
	. xy ( \ii1982|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \rstn_r_reg|qx_net  ),
	. f0 ( \io_phone_rst_inst|f_id[0]_net  )
);
defparam ii1982.PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.lut_0";
defparam ii1982.PCK_LOCATION = "C16R13.lp0.lut_0";
defparam ii1982.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii2082 (
	. xy ( \ii2082|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[11]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2082.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2082.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2082.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii1983 (
	. xy ( \ii1983|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  )
);
defparam ii1983.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.lut_0";
defparam ii1983.PCK_LOCATION = "C18R4.lp0.lut_0";
defparam ii1983.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
LUT6 ii2083 (
	. xy ( \ii2083|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[12]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2083.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2083.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2083.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28]|qx_net  ),
	. di ( \ii2176|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28] .always_en = 0;
LUT6 ii1984 (
	. xy ( \ii1984|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \mcu_arbiter_func_reg[0]|qx_net  ),
	. f1 ( \u_8051_u_h6_8051|port0o[0]_net  ),
	. f0 ( \ii1982_dup|xy_net  )
);
defparam ii1984.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii1984.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii1984.config_data = 64'b1000000010000000100000001000000010000000100000001000000010000000;
LUT6 ii2084 (
	. xy ( \ii2084|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[13]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2084.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2084.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2084.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]|qx_net  ),
	. di ( \ii2558|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .PLACE_LOCATION = "C20R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .PCK_LOCATION = "C20R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11] .always_en = 1;
LUT6 ii1985 (
	. xy ( \ii1985|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg|qx_net  ),
	. f1 ( \mipi_inst_u_mipi2|host_tx_payload_en_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii1985.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii1985.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii1985.config_data = 64'b0111111101111111011111110111111101111111011111110111111101111111;
LUT6 ii2085 (
	. xy ( \ii2085|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[14]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2085.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2085.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2085.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[25]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[25]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[25] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .PCK_LOCATION = "C20R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[0] .always_en = 1;
LUT6 ii2086 (
	. xy ( \ii2086|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[15]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2086.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2086.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2086.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7]|qx_net  ),
	. di ( \ii2518|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .PLACE_LOCATION = "C20R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .PCK_LOCATION = "C20R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[15] .always_en = 1;
LUT6 ii1987 (
	. xy ( \ii1987|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_fifo_vs_reg|qx_net  ),
	. f0 ( \ii1982_dup|xy_net  )
);
defparam ii1987.PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.lut_0";
defparam ii1987.PCK_LOCATION = "C16R15.lp0.lut_0";
defparam ii1987.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii2087 (
	. xy ( \ii2087|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[16]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2087.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2087.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2087.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11]|qx_net  ),
	. di ( \ii2369|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2341|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11] .always_en = 0;
LUT6 ii1988 (
	. xy ( \ii1988|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t85_out1_reg|qx_net  )
);
defparam ii1988.PLACE_LOCATION = "C6R25.le_tile.le_guts.lp0.lut_0";
defparam ii1988.PCK_LOCATION = "C6R25.lp0.lut_0";
defparam ii1988.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 ii2088 (
	. xy ( \ii2088|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[17]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2088.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2088.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2088.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .PCK_LOCATION = "C20R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[4] .always_en = 1;
LUT6 ii1989 (
	. xy ( \ii1989|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \glue_rx_packet_tx_packet_sc1_fifo_readen_reg|qx_net  )
);
defparam ii1989.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.lut_0";
defparam ii1989.PCK_LOCATION = "C14R7.lp0.lut_0";
defparam ii1989.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 ii1990 (
	. xy ( \ii1990|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg|qx_net  )
);
defparam ii1990.PLACE_LOCATION = "C14R6.le_tile.le_guts.lp0.lut_0";
defparam ii1990.PCK_LOCATION = "C14R6.lp0.lut_0";
defparam ii1990.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 ii2089 (
	. xy ( \ii2089|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[18]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2089.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2089.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2089.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2090 (
	. xy ( \ii2090|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[19]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2090.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2090.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2090.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2100 (
	. xy ( \ii2100|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[28]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[28]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2100.PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.lut_0";
defparam ii2100.PCK_LOCATION = "C14R27.lp0.lut_0";
defparam ii2100.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii1991 (
	. xy ( \ii1991|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0]|qx_net  )
);
defparam ii1991.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.lut_0";
defparam ii1991.PCK_LOCATION = "C20R23.lp0.lut_0";
defparam ii1991.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2091 (
	. xy ( \ii2091|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[1]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[1]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2091.PLACE_LOCATION = "C14R26.le_tile.le_guts.lp0.lut_0";
defparam ii2091.PCK_LOCATION = "C14R26.lp0.lut_0";
defparam ii2091.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2101 (
	. xy ( \ii2101|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[29]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[29]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2101.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2101.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2101.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8]|qx_net  ),
	. di ( \ii3108|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In2p_reg[8] .always_en = 1;
LUT6 ii1992 (
	. xy ( \ii1992|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10]|qx_net  )
);
defparam ii1992.PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.lut_0";
defparam ii1992.PCK_LOCATION = "C20R25.lp0.lut_0";
defparam ii1992.config_data = 64'b1110000011100000111000001110000011100000111000001110000011100000;
LUT6 ii2092 (
	. xy ( \ii2092|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[20]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2092.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2092.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2092.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2102 (
	. xy ( \ii2102|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[2]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[2]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2102.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2102.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2102.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg|qx_net  ),
	. di ( \ii3315|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_thd_vs_delay_flag_reg.always_en = 1;
LUT6 ii1993 (
	. xy ( \ii1993|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1]|qx_net  )
);
defparam ii1993.PLACE_LOCATION = "C18R24.le_tile.le_guts.lp0.lut_0";
defparam ii1993.PCK_LOCATION = "C18R24.lp0.lut_0";
defparam ii1993.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2093 (
	. xy ( \ii2093|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[21]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2093.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2093.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2093.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2103 (
	. xy ( \ii2103|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[30]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[30]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2103.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2103.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2103.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30]|qx_net  ),
	. di ( \ii2179|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29]|qx_net  ),
	. di ( \ii2177|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29] .always_en = 0;
LUT6 ii1994 (
	. xy ( \ii1994|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2]|qx_net  )
);
defparam ii1994.PLACE_LOCATION = "C18R24.le_tile.le_guts.lp0.lut_0";
defparam ii1994.PCK_LOCATION = "C18R24.lp0.lut_0";
defparam ii1994.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2094 (
	. xy ( \ii2094|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[22]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2094.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2094.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2094.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2104 (
	. xy ( \ii2104|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[31]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[31]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2104.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2104.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2104.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii1995 (
	. xy ( \ii1995|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3]|qx_net  )
);
defparam ii1995.PLACE_LOCATION = "C18R24.le_tile.le_guts.lp0.lut_0";
defparam ii1995.PCK_LOCATION = "C18R24.lp0.lut_0";
defparam ii1995.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2095 (
	. xy ( \ii2095|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[23]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2095.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2095.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2095.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2105 (
	. xy ( \ii2105|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[3]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[3]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2105.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2105.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2105.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[26]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[26]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[26] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .PCK_LOCATION = "C20R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[1] .always_en = 1;
LUT6 ii1996 (
	. xy ( \ii1996|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4]|qx_net  )
);
defparam ii1996.PLACE_LOCATION = "C18R24.le_tile.le_guts.lp0.lut_0";
defparam ii1996.PCK_LOCATION = "C18R24.lp0.lut_0";
defparam ii1996.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2096 (
	. xy ( \ii2096|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[24]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2096.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2096.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2096.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2106 (
	. xy ( \ii2106|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[4]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[4]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2106.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2106.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2106.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[16] .always_en = 1;
LUT6 ii1997 (
	. xy ( \ii1997|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5]|qx_net  )
);
defparam ii1997.PLACE_LOCATION = "C18R24.le_tile.le_guts.lp0.lut_0";
defparam ii1997.PCK_LOCATION = "C18R24.lp0.lut_0";
defparam ii1997.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2097 (
	. xy ( \ii2097|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[25]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2097.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2097.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2097.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2107 (
	. xy ( \ii2107|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[5]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[5]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2107.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2107.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2107.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii1998 (
	. xy ( \ii1998|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6]|qx_net  )
);
defparam ii1998.PLACE_LOCATION = "C18R24.le_tile.le_guts.lp0.lut_0";
defparam ii1998.PCK_LOCATION = "C18R24.lp0.lut_0";
defparam ii1998.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2098 (
	. xy ( \ii2098|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[26]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[26]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2098.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2098.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2098.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2108 (
	. xy ( \ii2108|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[6]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[6]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2108.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2108.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2108.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .PCK_LOCATION = "C20R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[5] .always_en = 1;
LUT6 ii1999 (
	. xy ( \ii1999|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t47_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7]|qx_net  )
);
defparam ii1999.PLACE_LOCATION = "C20R24.le_tile.le_guts.lp0.lut_0";
defparam ii1999.PCK_LOCATION = "C20R24.lp0.lut_0";
defparam ii1999.config_data = 64'b1010110010101100101011001010110010101100101011001010110010101100;
LUT6 ii2099 (
	. xy ( \ii2099|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[27]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[27]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2099.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2099.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2099.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2109 (
	. xy ( \ii2109|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[7]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[7]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2109.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2109.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2109.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2110 (
	. xy ( \ii2110|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[8]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[8]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2110.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2110.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2110.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2111 (
	. xy ( \ii2111|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[9]|qx_net  ),
	. f1 ( \mcu_arbiter_u_pfifo_u_inst|dout[9]_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2111.PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.lut_0";
defparam ii2111.PCK_LOCATION = "C14R28.lp0.lut_0";
defparam ii2111.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2112 (
	. xy ( \ii2112|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_mipi_sel_reg|qx_net  ),
	. f0 ( \ii2050|xy_net  )
);
defparam ii2112.PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.lut_0";
defparam ii2112.PCK_LOCATION = "C10R15.lp0.lut_0";
defparam ii2112.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG glue_rx_packet_tx_packet_sc_vs_reg (
	. qx ( \glue_rx_packet_tx_packet_sc_vs_reg|qx_net  ),
	. di ( \ii2141|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_sc_vs_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.init = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc_vs_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_sc_vs_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.PCK_LOCATION = "C20R18.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc_vs_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_sc_vs_reg.always_en = 1;
LUT6 ii2113 (
	. xy ( \ii2113|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_fifo_readen_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  )
);
defparam ii2113.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2113.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2113.config_data = 64'b1110111011101110111011101110111011101110111011101110111011101110;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31]|qx_net  ),
	. di ( \ii2180|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .PCK_LOCATION = "C14R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0] .always_en = 1;
LUT6 ii2114 (
	. xy ( \ii2114|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_memack_reg|qx_net  ),
	. f4 ( \mcu_arbiter_u_emif2apb_memack_reg|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_memack_reg|qx_net  ),
	. f1 ( \mcu_arbiter_data_sel_reg|qx_net  ),
	. f0 ( \mcu_arbiter_apb_sel_reg|qx_net  )
);
defparam ii2114.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.lut_0";
defparam ii2114.PCK_LOCATION = "C4R18.lp0.lut_0";
defparam ii2114.config_data = 64'b1111000011101110111100000100010011110000101010101111000000000000;
LUT6 ii2115 (
	. xy ( \ii2115|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[8]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[24]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[16]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[0]_net  )
);
defparam ii2115.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2115.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2115.config_data = 64'b1111000011110000110011001100110011111111000000001010101010101010;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[27]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[27]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[27] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .PCK_LOCATION = "C20R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[2] .always_en = 1;
LUT6 ii2116 (
	. xy ( \ii2116|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[0]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2115|xy_net  )
);
defparam ii2116.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2116.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2116.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .PCK_LOCATION = "C4R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[17] .always_en = 1;
LUT6 ii2117 (
	. xy ( \ii2117|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[9]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[25]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[1]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[17]_net  )
);
defparam ii2117.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2117.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2117.config_data = 64'b1111000011110000101010101010101011111111000000001100110011001100;
LUT6 ii2118 (
	. xy ( \ii2118|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[1]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[1]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2117|xy_net  )
);
defparam ii2118.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2118.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2118.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .PCK_LOCATION = "C20R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[6] .always_en = 1;
LUT6 ii2119 (
	. xy ( \ii2119|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[2]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[26]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[18]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[10]_net  )
);
defparam ii2119.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2119.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2119.config_data = 64'b1111000011110000110011001100110010101010101010101111111100000000;
LUT6 ii2120 (
	. xy ( \ii2120|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[2]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[2]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2119|xy_net  )
);
defparam ii2120.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2120.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2120.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
LUT6 ii2121 (
	. xy ( \ii2121|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[3]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[27]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[19]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[11]_net  )
);
defparam ii2121.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2121.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2121.config_data = 64'b1111000011110000110011001100110010101010101010101111111100000000;
LUT6 ii2122 (
	. xy ( \ii2122|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[3]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[3]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2121|xy_net  )
);
defparam ii2122.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2122.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2122.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
LUT6 ii2123 (
	. xy ( \ii2123|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[4]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[28]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[20]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[12]_net  )
);
defparam ii2123.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2123.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2123.config_data = 64'b1111000011110000110011001100110010101010101010101111111100000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32]|qx_net  ),
	. di ( \ii2181|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32] .always_en = 0;
ADD1_A carry_12_2__ADD_10 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10]|qx_net  ),
	. ci ( \carry_12_2__ADD_9|co_net  ),
	. co ( \carry_12_2__ADD_10|co_net  ),
	. s ( \carry_12_2__ADD_10|s_net  )
);
defparam carry_12_2__ADD_10.PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_10.a_inv = "false";
defparam carry_12_2__ADD_10.PCK_LOCATION = "C16R5.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0]|qx_net  ),
	. di ( \ii2608|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1] .always_en = 1;
SPRAM_2Kx32 glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram (
	. clk ( \u_pll_pll_u0|CO0_net  ),
	. addr ( {
		/* addr [10] */ \ii1992|xy_net ,
		/* addr [9] */ \ii2001|xy_net ,
		/* addr [8] */ \ii2000|xy_net ,
		/* addr [7] */ \ii1999|xy_net ,
		/* addr [6] */ \ii1998|xy_net ,
		/* addr [5] */ \ii1997|xy_net ,
		/* addr [4] */ \ii1996|xy_net ,
		/* addr [3] */ \ii1995|xy_net ,
		/* addr [2] */ \ii1994|xy_net ,
		/* addr [1] */ \ii1993|xy_net ,
		/* addr [0] */ \ii1991|xy_net 
	} ),
	. datai ( {
		/* datai [31] */ \GND_0_inst|Y_net ,
		/* datai [30] */ \GND_0_inst|Y_net ,
		/* datai [29] */ \GND_0_inst|Y_net ,
		/* datai [28] */ \GND_0_inst|Y_net ,
		/* datai [27] */ \GND_0_inst|Y_net ,
		/* datai [26] */ \GND_0_inst|Y_net ,
		/* datai [25] */ \GND_0_inst|Y_net ,
		/* datai [24] */ \GND_0_inst|Y_net ,
		/* datai [23] */ \GND_0_inst|Y_net ,
		/* datai [22] */ \GND_0_inst|Y_net ,
		/* datai [21] */ \GND_0_inst|Y_net ,
		/* datai [20] */ \GND_0_inst|Y_net ,
		/* datai [19] */ \GND_0_inst|Y_net ,
		/* datai [18] */ \GND_0_inst|Y_net ,
		/* datai [17] */ \GND_0_inst|Y_net ,
		/* datai [16] */ \GND_0_inst|Y_net ,
		/* datai [15] */ \GND_0_inst|Y_net ,
		/* datai [14] */ \GND_0_inst|Y_net ,
		/* datai [13] */ \GND_0_inst|Y_net ,
		/* datai [12] */ \GND_0_inst|Y_net ,
		/* datai [11] */ \GND_0_inst|Y_net ,
		/* datai [10] */ \GND_0_inst|Y_net ,
		/* datai [9] */ \GND_0_inst|Y_net ,
		/* datai [8] */ \GND_0_inst|Y_net ,
		/* datai [7] */ \GND_0_inst|Y_net ,
		/* datai [6] */ \GND_0_inst|Y_net ,
		/* datai [5] */ \GND_0_inst|Y_net ,
		/* datai [4] */ \GND_0_inst|Y_net ,
		/* datai [3] */ \GND_0_inst|Y_net ,
		/* datai [2] */ \GND_0_inst|Y_net ,
		/* datai [1] */ \GND_0_inst|Y_net ,
		/* datai [0] */ \GND_0_inst|Y_net 
	} ),
	. ceb ( \GND_0_inst|Y_net  ),
	. web ( \VCC_0_inst|Y_net  ),
	. datao ( {
		/* datao [31] (nc) */ nc460 ,
		/* datao [30] (nc) */ nc461 ,
		/* datao [29] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[29]_net ,
		/* datao [28] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[28]_net ,
		/* datao [27] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[27]_net ,
		/* datao [26] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[26]_net ,
		/* datao [25] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[25]_net ,
		/* datao [24] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[24]_net ,
		/* datao [23] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[23]_net ,
		/* datao [22] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[22]_net ,
		/* datao [21] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[21]_net ,
		/* datao [20] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[20]_net ,
		/* datao [19] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[19]_net ,
		/* datao [18] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[18]_net ,
		/* datao [17] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[17]_net ,
		/* datao [16] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[16]_net ,
		/* datao [15] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[15]_net ,
		/* datao [14] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[14]_net ,
		/* datao [13] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[13]_net ,
		/* datao [12] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[12]_net ,
		/* datao [11] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[11]_net ,
		/* datao [10] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[10]_net ,
		/* datao [9] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[9]_net ,
		/* datao [8] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[8]_net ,
		/* datao [7] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[7]_net ,
		/* datao [6] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[6]_net ,
		/* datao [5] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[5]_net ,
		/* datao [4] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[4]_net ,
		/* datao [3] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[3]_net ,
		/* datao [2] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[2]_net ,
		/* datao [1] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[1]_net ,
		/* datao [0] */ \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[0]_net 
	} )
);
defparam glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram.PLACE_LOCATION = "C23R29.spram_2kx32_wrap0.spram_2kx32";
defparam glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram.PCK_LOCATION = "NONE";
defparam glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram.init_file = "src/emb_2160_1080_to_1440_720.dat";
LUT6 ii2124 (
	. xy ( \ii2124|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[4]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[4]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2123|xy_net  )
);
defparam ii2124.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2124.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2124.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
ADD1_A carry_12_2__ADD_11 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11]|qx_net  ),
	. ci ( \carry_12_2__ADD_10|co_net  ),
	. co ( ),
	. s ( \carry_12_2__ADD_11|s_net  )
);
defparam carry_12_2__ADD_11.PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_2__ADD_11.a_inv = "false";
defparam carry_12_2__ADD_11.PCK_LOCATION = "C16R5.lp0.add2.add0";
LUT6 ii2125 (
	. xy ( \ii2125|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[5]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[29]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[21]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[13]_net  )
);
defparam ii2125.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2125.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2125.config_data = 64'b1111000011110000110011001100110010101010101010101111111100000000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[28]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[28]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[3] .always_en = 1;
LUT6 ii2126 (
	. xy ( \ii2126|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[5]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[5]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2125|xy_net  )
);
defparam ii2126.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2126.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2126.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[18] .always_en = 1;
LUT6 ii2127 (
	. xy ( \ii2127|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[6]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[30]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[22]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[14]_net  )
);
defparam ii2127.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2127.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2127.config_data = 64'b1111000011110000110011001100110010101010101010101111111100000000;
LUT6 ii2128 (
	. xy ( \ii2128|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[6]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[6]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2127|xy_net  )
);
defparam ii2128.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2128.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2128.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .PCK_LOCATION = "C20R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In3p_reg[7] .always_en = 1;
LUT6 ii2129 (
	. xy ( \ii2129|xy_net  ),
	. f5 ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. f4 ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. f3 ( \mcu_arbiter_u_psram_u_psram|datao[7]_net  ),
	. f2 ( \mcu_arbiter_u_psram_u_psram|datao[31]_net  ),
	. f1 ( \mcu_arbiter_u_psram_u_psram|datao[23]_net  ),
	. f0 ( \mcu_arbiter_u_psram_u_psram|datao[15]_net  )
);
defparam ii2129.PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.lut_0";
defparam ii2129.PCK_LOCATION = "C18R27.lp0.lut_0";
defparam ii2129.config_data = 64'b1111000011110000110011001100110010101010101010101111111100000000;
LUT6 ii2130 (
	. xy ( \ii2130|xy_net  ),
	. f5 ( ),
	. f4 ( \mcu_arbiter_u_emif2apb_memdatai_reg[7]|qx_net  ),
	. f3 ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. f2 ( \mcu_arbiter_reg_din_reg[7]|qx_net  ),
	. f1 ( \mcu_arbiter_apb_sel_reg|qx_net  ),
	. f0 ( \ii2129|xy_net  )
);
defparam ii2130.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.lut_0";
defparam ii2130.PCK_LOCATION = "C4R20.lp0.lut_0";
defparam ii2130.config_data = 64'b1111000011101110111100000010001011110000111011101111000000100010;
LUT6 ii2131 (
	. xy ( \ii2131|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mcu_arbiter_u_psram_memack_reg|qx_net  ),
	. f0 ( \mcu_arbiter_code_sel_reg|qx_net  )
);
defparam ii2131.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.lut_0";
defparam ii2131.PCK_LOCATION = "C4R18.lp0.lut_0";
defparam ii2131.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii2132 (
	. xy ( \ii2132|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \mipi_inst_u_mipi_pll|LOCK_net  ),
	. f1 ( \mipi_inst_u_mipi2|tx_dphy_rdy_net  ),
	. f0 ( \mipi_inst_u_mipi1|tx_dphy_rdy_net  )
);
defparam ii2132.PLACE_LOCATION = "C6R11.le_tile.le_guts.lp0.lut_0";
defparam ii2132.PCK_LOCATION = "C6R11.lp0.lut_0";
defparam ii2132.config_data = 64'b1000000010000000100000001000000010000000100000001000000010000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33]|qx_net  ),
	. di ( \ii2182|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .PCK_LOCATION = "C20R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t46_reg_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_10__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .PCK_LOCATION = "C18R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[0] .always_en = 1;
LUT6 ii2134 (
	. xy ( \ii2134|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. f2 ( \glue_pasm_cmd_rq_o_reg|qx_net  ),
	. f1 ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2134.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.lut_0";
defparam ii2134.PCK_LOCATION = "C14R30.lp0.lut_0";
defparam ii2134.config_data = 64'b1011101110110000101110111011000010111011101100001011101110110000;
LUT6 ii2135 (
	. xy ( \ii2135|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rd_cmd_flag_d_reg|qx_net  ),
	. f3 ( \glue_pasm_tx_act_d_reg|qx_net  ),
	. f2 ( \glue_pasm_packet_finish_reg|qx_net  ),
	. f1 ( \mipi_inst_u_mipi2|host_tx_active_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2135.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2135.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2135.config_data = 64'b0000000000000000111110111111000000000000000000001111101111110000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[29]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[29]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[29] .always_en = 1;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[30]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[30]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[30] .always_en = 1;
ADD1_A carry_9_8__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_8__ADD_0|co_net  ),
	. s ( \carry_9_8__ADD_0|s_net  )
);
defparam carry_9_8__ADD_0.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_0.a_inv = "true";
defparam carry_9_8__ADD_0.PCK_LOCATION = "C18R9.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[4] .always_en = 1;
LUT6 ii2136 (
	. xy ( \ii2136|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mipi_inst_u_mipi2|host_tx_active_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2136.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.lut_0";
defparam ii2136.PCK_LOCATION = "C14R30.lp0.lut_0";
defparam ii2136.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[4]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf.PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf.PCK_LOCATION = "C14R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .PLACE_LOCATION = "C6R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .PCK_LOCATION = "C6R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[3] .always_en = 1;
ADD1_A carry_9_8__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1]|qx_net  ),
	. ci ( \carry_9_8__ADD_0|co_net  ),
	. co ( \carry_9_8__ADD_1|co_net  ),
	. s ( \carry_9_8__ADD_1|s_net  )
);
defparam carry_9_8__ADD_1.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_1.a_inv = "true";
defparam carry_9_8__ADD_1.PCK_LOCATION = "C18R9.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[20] .always_en = 1;
LUT6 ii2137 (
	. xy ( \ii2137|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rd_start_s_reg|qx_net  ),
	. f0 ( \glue_rd_start_d_reg|qx_net  )
);
defparam ii2137.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii2137.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii2137.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg|qx_net  ),
	. di ( \ii2292|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.PCK_LOCATION = "C14R25.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg.always_en = 1;
ADD1_A carry_9_8__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2]|qx_net  ),
	. ci ( \carry_9_8__ADD_1|co_net  ),
	. co ( \carry_9_8__ADD_2|co_net  ),
	. s ( \carry_9_8__ADD_2|s_net  )
);
defparam carry_9_8__ADD_2.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_2.a_inv = "true";
defparam carry_9_8__ADD_2.PCK_LOCATION = "C18R9.lp0.add2.add0";
LUT6 ii2138 (
	. xy ( \ii2138|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \mcu_arbiter_func_reg[0]|qx_net  ),
	. f1 ( \u_8051_u_h6_8051|port0o[1]_net  ),
	. f0 ( \ii1982_dup|xy_net  )
);
defparam ii2138.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii2138.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii2138.config_data = 64'b1000000010000000100000001000000010000000100000001000000010000000;
REG glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg (
	. qx ( \glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg|qx_net  ),
	. di ( \ii2380|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.init = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.PLACE_LOCATION = "C10R6.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.PCK_LOCATION = "C10R6.lp0.reg0";
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg.always_en = 1;
FIFO18K glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst (
	. dout ( {
		/* dout [63] (nc) */ nc462 ,
		/* dout [62] (nc) */ nc463 ,
		/* dout [61] (nc) */ nc464 ,
		/* dout [60] (nc) */ nc465 ,
		/* dout [59] (nc) */ nc466 ,
		/* dout [58] (nc) */ nc467 ,
		/* dout [57] (nc) */ nc468 ,
		/* dout [56] (nc) */ nc469 ,
		/* dout [55] (nc) */ nc470 ,
		/* dout [54] (nc) */ nc471 ,
		/* dout [53] (nc) */ nc472 ,
		/* dout [52] (nc) */ nc473 ,
		/* dout [51] (nc) */ nc474 ,
		/* dout [50] (nc) */ nc475 ,
		/* dout [49] (nc) */ nc476 ,
		/* dout [48] (nc) */ nc477 ,
		/* dout [47] (nc) */ nc478 ,
		/* dout [46] (nc) */ nc479 ,
		/* dout [45] (nc) */ nc480 ,
		/* dout [44] (nc) */ nc481 ,
		/* dout [43] (nc) */ nc482 ,
		/* dout [42] (nc) */ nc483 ,
		/* dout [41] (nc) */ nc484 ,
		/* dout [40] (nc) */ nc485 ,
		/* dout [39] (nc) */ nc486 ,
		/* dout [38] (nc) */ nc487 ,
		/* dout [37] (nc) */ nc488 ,
		/* dout [36] (nc) */ nc489 ,
		/* dout [35] (nc) */ nc490 ,
		/* dout [34] (nc) */ nc491 ,
		/* dout [33] (nc) */ nc492 ,
		/* dout [32] (nc) */ nc493 ,
		/* dout [31] (nc) */ nc494 ,
		/* dout [30] (nc) */ nc495 ,
		/* dout [29] (nc) */ nc496 ,
		/* dout [28] (nc) */ nc497 ,
		/* dout [27] (nc) */ nc498 ,
		/* dout [26] (nc) */ nc499 ,
		/* dout [25] (nc) */ nc500 ,
		/* dout [24] (nc) */ nc501 ,
		/* dout [23] (nc) */ nc502 ,
		/* dout [22] (nc) */ nc503 ,
		/* dout [21] (nc) */ nc504 ,
		/* dout [20] (nc) */ nc505 ,
		/* dout [19] (nc) */ nc506 ,
		/* dout [18] (nc) */ nc507 ,
		/* dout [17] (nc) */ nc508 ,
		/* dout [16] (nc) */ nc509 ,
		/* dout [15] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[15]_net ,
		/* dout [14] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[14]_net ,
		/* dout [13] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[13]_net ,
		/* dout [12] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[12]_net ,
		/* dout [11] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[11]_net ,
		/* dout [10] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[10]_net ,
		/* dout [9] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[9]_net ,
		/* dout [8] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[8]_net ,
		/* dout [7] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[7]_net ,
		/* dout [6] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[6]_net ,
		/* dout [5] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[5]_net ,
		/* dout [4] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[4]_net ,
		/* dout [3] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[3]_net ,
		/* dout [2] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[2]_net ,
		/* dout [1] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[1]_net ,
		/* dout [0] */ \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[0]_net 
	} ),
	. doutp ( )
,
	. din ( {
		/* din [63] */ \GND_0_inst|Y_net ,
		/* din [62] */ \GND_0_inst|Y_net ,
		/* din [61] */ \GND_0_inst|Y_net ,
		/* din [60] */ \GND_0_inst|Y_net ,
		/* din [59] */ \GND_0_inst|Y_net ,
		/* din [58] */ \GND_0_inst|Y_net ,
		/* din [57] */ \GND_0_inst|Y_net ,
		/* din [56] */ \GND_0_inst|Y_net ,
		/* din [55] */ \GND_0_inst|Y_net ,
		/* din [54] */ \GND_0_inst|Y_net ,
		/* din [53] */ \GND_0_inst|Y_net ,
		/* din [52] */ \GND_0_inst|Y_net ,
		/* din [51] */ \GND_0_inst|Y_net ,
		/* din [50] */ \GND_0_inst|Y_net ,
		/* din [49] */ \GND_0_inst|Y_net ,
		/* din [48] */ \GND_0_inst|Y_net ,
		/* din [47] */ \GND_0_inst|Y_net ,
		/* din [46] */ \GND_0_inst|Y_net ,
		/* din [45] */ \GND_0_inst|Y_net ,
		/* din [44] */ \GND_0_inst|Y_net ,
		/* din [43] */ \GND_0_inst|Y_net ,
		/* din [42] */ \GND_0_inst|Y_net ,
		/* din [41] */ \GND_0_inst|Y_net ,
		/* din [40] */ \GND_0_inst|Y_net ,
		/* din [39] */ \GND_0_inst|Y_net ,
		/* din [38] */ \GND_0_inst|Y_net ,
		/* din [37] */ \GND_0_inst|Y_net ,
		/* din [36] */ \GND_0_inst|Y_net ,
		/* din [35] */ \GND_0_inst|Y_net ,
		/* din [34] */ \GND_0_inst|Y_net ,
		/* din [33] */ \GND_0_inst|Y_net ,
		/* din [32] */ \GND_0_inst|Y_net ,
		/* din [31] */ \GND_0_inst|Y_net ,
		/* din [30] */ \GND_0_inst|Y_net ,
		/* din [29] */ \GND_0_inst|Y_net ,
		/* din [28] */ \GND_0_inst|Y_net ,
		/* din [27] */ \GND_0_inst|Y_net ,
		/* din [26] */ \GND_0_inst|Y_net ,
		/* din [25] */ \GND_0_inst|Y_net ,
		/* din [24] */ \GND_0_inst|Y_net ,
		/* din [23] */ \GND_0_inst|Y_net ,
		/* din [22] */ \GND_0_inst|Y_net ,
		/* din [21] */ \GND_0_inst|Y_net ,
		/* din [20] */ \GND_0_inst|Y_net ,
		/* din [19] */ \GND_0_inst|Y_net ,
		/* din [18] */ \GND_0_inst|Y_net ,
		/* din [17] */ \GND_0_inst|Y_net ,
		/* din [16] */ \GND_0_inst|Y_net ,
		/* din [15] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[23]|qx_net ,
		/* din [14] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[22]|qx_net ,
		/* din [13] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[21]|qx_net ,
		/* din [12] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[20]|qx_net ,
		/* din [11] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[19]|qx_net ,
		/* din [10] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18]|qx_net ,
		/* din [9] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17]|qx_net ,
		/* din [8] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16]|qx_net ,
		/* din [7] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[31]|qx_net ,
		/* din [6] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[30]|qx_net ,
		/* din [5] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[29]|qx_net ,
		/* din [4] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[28]|qx_net ,
		/* din [3] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[27]|qx_net ,
		/* din [2] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[26]|qx_net ,
		/* din [1] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[25]|qx_net ,
		/* din [0] */ \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[24]|qx_net 
	} ),
	. dinp ( {
		/* dinp [7] */ \GND_0_inst|Y_net ,
		/* dinp [6] */ \GND_0_inst|Y_net ,
		/* dinp [5] */ \GND_0_inst|Y_net ,
		/* dinp [4] */ \GND_0_inst|Y_net ,
		/* dinp [3] */ \GND_0_inst|Y_net ,
		/* dinp [2] */ \GND_0_inst|Y_net ,
		/* dinp [1] */ \GND_0_inst|Y_net ,
		/* dinp [0] */ \GND_0_inst|Y_net 
	} ),
	. writeclk ( \u_pll_pll_u0|CO0_net  ),
	. readclk ( \u_gbuf_u_gbuf|out_net  ),
	. writeen ( \ii1988|xy_net  ),
	. readen ( \ii1985|xy_net  ),
	. reset ( \ii1987|xy_net  ),
	. regce ( \VCC_0_inst|Y_net  ),
	. writesave ( \GND_0_inst|Y_net  ),
	. writedrop ( \GND_0_inst|Y_net  ),
	. full ( ),
	. empty ( ),
	. almostfull ( ),
	. almostempty ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|almostempty_net  ),
	. overflow ( ),
	. underflow ( ),
	. eccoutdberr ( ),
	. eccoutsberr ( ),
	. eccreadaddr ( )
,
	. eccindberr ( \GND_0_inst|Y_net  ),
	. eccinsberr ( \GND_0_inst|Y_net  ),
	. writedropflag ( )
);
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.eccwriteen = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.writeclk_inv = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.eccreaden = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.readclk_inv = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.use_parity = 0;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.outreg = 1;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.almostfullth = 988;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.almostemptyth = 512;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.writewidth = 18;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.readwidth = 18;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.peek = 1;
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.PLACE_LOCATION = "C12R21.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst.PCK_LOCATION = "C12R21.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
ADD1_A carry_9_8__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3]|qx_net  ),
	. ci ( \carry_9_8__ADD_2|co_net  ),
	. co ( \carry_9_8__ADD_3|co_net  ),
	. s ( \carry_9_8__ADD_3|s_net  )
);
defparam carry_9_8__ADD_3.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_3.a_inv = "true";
defparam carry_9_8__ADD_3.PCK_LOCATION = "C18R9.lp0.add2.add0";
LUT6 ii2139 (
	. xy ( \ii2139|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|almostempty_net  ),
	. f0 ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|almostempty_net  )
);
defparam ii2139.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2139.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2139.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii2140 (
	. xy ( \ii2140|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|empty_net  )
);
defparam ii2140.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam ii2140.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam ii2140.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
ADD1_A carry_9_8__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4]|qx_net  ),
	. ci ( \carry_9_8__ADD_3|co_net  ),
	. co ( \carry_9_8__ADD_4|co_net  ),
	. s ( \carry_9_8__ADD_4|s_net  )
);
defparam carry_9_8__ADD_4.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_4.a_inv = "true";
defparam carry_9_8__ADD_4.PCK_LOCATION = "C18R9.lp0.add2.add0";
LUT6 ii2141 (
	. xy ( \ii2141|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rstsf_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rstsf_reg[0]|qx_net  )
);
defparam ii2141.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii2141.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii2141.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
ADD1_A carry_9_8__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5]|qx_net  ),
	. ci ( \carry_9_8__ADD_4|co_net  ),
	. co ( \carry_9_8__ADD_5|co_net  ),
	. s ( \carry_9_8__ADD_5|s_net  )
);
defparam carry_9_8__ADD_5.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_5.a_inv = "true";
defparam carry_9_8__ADD_5.PCK_LOCATION = "C18R9.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. di ( \ii2613|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .PCK_LOCATION = "C16R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0] .always_en = 1;
LUT6 ii2142 (
	. xy ( \ii2142|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \ii2141|xy_net  )
);
defparam ii2142.PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.lut_0";
defparam ii2142.PCK_LOCATION = "C20R13.lp0.lut_0";
defparam ii2142.config_data = 64'b0101010101010101010101010101010101010101010101010101010101010101;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[27]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf.PLACE_LOCATION = "C4R12.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf.PCK_LOCATION = "C4R12.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
ADD1_A carry_9_8__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6]|qx_net  ),
	. ci ( \carry_9_8__ADD_5|co_net  ),
	. co ( \carry_9_8__ADD_6|co_net  ),
	. s ( \carry_9_8__ADD_6|s_net  )
);
defparam carry_9_8__ADD_6.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_6.a_inv = "true";
defparam carry_9_8__ADD_6.PCK_LOCATION = "C18R9.lp0.add2.add0";
LUT6 ii2143 (
	. xy ( \ii2143|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]|qx_net  )
);
defparam ii2143.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2143.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2143.config_data = 64'b0100000000000000000000000000000000000000000000000000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34]|qx_net  ),
	. di ( \ii2183|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34] .always_en = 0;
ADD1_A carry_9_8__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7]|qx_net  ),
	. ci ( \carry_9_8__ADD_6|co_net  ),
	. co ( \carry_9_8__ADD_7|co_net  ),
	. s ( \carry_9_8__ADD_7|s_net  )
);
defparam carry_9_8__ADD_7.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_7.a_inv = "true";
defparam carry_9_8__ADD_7.PCK_LOCATION = "C18R9.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .PLACE_LOCATION = "C20R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .PCK_LOCATION = "C20R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_10__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .PCK_LOCATION = "C18R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[1] .always_en = 1;
LUT6 ii2144 (
	. xy ( \ii2144|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg|qx_net  ),
	. f3 ( \mipi_inst_u_mipi2|host_tx_payload_en_last_net  ),
	. f2 ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. f1 ( \ii2143|xy_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2144.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2144.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2144.config_data = 64'b1101010111111111100000001000000001010101111111110000000000000000;
ADD1_A carry_9_8__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_8__ADD_7|co_net  ),
	. co ( \carry_9_8__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_8__ADD_8.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_8__ADD_8.a_inv = "false";
defparam carry_9_8__ADD_8.PCK_LOCATION = "C18R10.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .PCK_LOCATION = "C10R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[0] .always_en = 1;
LUT6 ii2145 (
	. xy ( \ii2145|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_req_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg|qx_net  ),
	. f2 ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. f1 ( \ii2143|xy_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2145.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.lut_0";
defparam ii2145.PCK_LOCATION = "C14R29.lp0.lut_0";
defparam ii2145.config_data = 64'b1101111111001100010111110000000011011111110011000101111100000000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[31]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[31]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[31] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .PCK_LOCATION = "C20R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_In1p_reg[5] .always_en = 1;
LUT6 ii2146 (
	. xy ( \ii2146|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  )
);
defparam ii2146.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2146.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2146.config_data = 64'b0000000010101110000000001010111000000000101011100000000010101110;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[4] .always_en = 1;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg|qx_net  ),
	. di ( \ii2144|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.PCK_LOCATION = "C14R29.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_packet_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[21] .always_en = 1;
LUT6 ii2147 (
	. xy ( \ii2147|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[10]|qx_net  )
);
defparam ii2147.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2147.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2147.config_data = 64'b1010101010101010101010101010101010101000000000000000000000000000;
LUT6 ii2148 (
	. xy ( \ii2148|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[11]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg|qx_net  ),
	. f0 ( \ii2147|xy_net  )
);
defparam ii2148.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2148.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2148.config_data = 64'b0000000000000000000000000000000000000000000000000101010100010000;
LUT6 ii2149 (
	. xy ( \ii2149|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2149.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.lut_0";
defparam ii2149.PCK_LOCATION = "C14R30.lp0.lut_0";
defparam ii2149.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
LUT6 ii2150 (
	. xy ( \ii2150|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  )
);
defparam ii2150.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2150.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2150.config_data = 64'b0100010001000100010001000100010001000100010001000100010001000100;
LUT6 ii2151 (
	. xy ( \ii2151|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2151.PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.lut_0";
defparam ii2151.PCK_LOCATION = "C14R19.lp0.lut_0";
defparam ii2151.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. di ( \ii2659|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1] .always_en = 1;
LUT6 ii2152 (
	. xy ( \ii2152|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  )
);
defparam ii2152.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2152.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2152.config_data = 64'b0000101100001011000010110000101100001011000010110000101100001011;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.PCK_LOCATION = "C14R22.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg.always_en = 1;
LUT6 ii2153 (
	. xy ( \ii2153|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  ),
	. f2 ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2153.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2153.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2153.config_data = 64'b1111111110110011101100111011001111111111101100111011001110110011;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35]|qx_net  ),
	. di ( \ii2184|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_10__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .PCK_LOCATION = "C18R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[2] .always_en = 1;
LUT6 ii2154 (
	. xy ( \ii2154|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2154.PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.lut_0";
defparam ii2154.PCK_LOCATION = "C14R19.lp0.lut_0";
defparam ii2154.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .PCK_LOCATION = "C10R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[1] .always_en = 1;
LUT6 ii2155 (
	. xy ( \ii2155|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2155.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2155.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2155.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2156 (
	. xy ( \ii2156|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2156.PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.lut_0";
defparam ii2156.PCK_LOCATION = "C14R19.lp0.lut_0";
defparam ii2156.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[22] .always_en = 1;
LUT6 ii2157 (
	. xy ( \ii2157|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2157.PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.lut_0";
defparam ii2157.PCK_LOCATION = "C14R19.lp0.lut_0";
defparam ii2157.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2158 (
	. xy ( \ii2158|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2158.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2158.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2158.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2159 (
	. xy ( \ii2159|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2159.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2159.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2159.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2160 (
	. xy ( \ii2160|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2160.PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.lut_0";
defparam ii2160.PCK_LOCATION = "C14R19.lp0.lut_0";
defparam ii2160.config_data = 64'b0101111101011100010111110101110001011111010111000101111101011100;
LUT6 ii2161 (
	. xy ( \ii2161|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[0]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2161.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2161.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2161.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0]|qx_net  ),
	. di ( \ii2584|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. di ( \ii2711|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2] .always_en = 1;
LUT6 ii2162 (
	. xy ( \ii2162|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[1]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2162.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2162.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2162.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2163 (
	. xy ( \ii2163|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[2]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2163.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2163.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2163.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36]|qx_net  ),
	. di ( \ii2185|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_10__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .PCK_LOCATION = "C18R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[3] .always_en = 1;
LUT6 ii2164 (
	. xy ( \ii2164|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[3]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2164.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2164.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2164.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .PCK_LOCATION = "C10R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[2] .always_en = 1;
LUT6 ii2165 (
	. xy ( \ii2165|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2165.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2165.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2165.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG mcu_arbiter_u_emif2apb_memack_reg (
	. qx ( \mcu_arbiter_u_emif2apb_memack_reg|qx_net  ),
	. di ( \ii3340|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_emif2apb_memack_reg.latch_mode = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.init = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.PLACE_LOCATION = "C4R17.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_memack_reg.sr_inv = 1;
defparam mcu_arbiter_u_emif2apb_memack_reg.sync_mode = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.no_sr = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.sr_value = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.PCK_LOCATION = "C4R17.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_memack_reg.clk_inv = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.en_inv = 0;
defparam mcu_arbiter_u_emif2apb_memack_reg.always_en = 1;
LUT6 ii2166 (
	. xy ( \ii2166|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2152|xy_net  )
);
defparam ii2166.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2166.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2166.config_data = 64'b1010001010100010101000101010001010100010101000101010001010100010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[23] .always_en = 1;
LUT6 ii2167 (
	. xy ( \ii2167|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_fifo_empty_reg|qx_net  )
);
defparam ii2167.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2167.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2167.config_data = 64'b0100000001000000010000000100000001000000010000000100000001000000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[17]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2168 (
	. xy ( \ii2168|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2168.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2168.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2168.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
LUT6 ii2169 (
	. xy ( \ii2169|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[5]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2169.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2169.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2169.config_data = 64'b1100110011001100010001001100000011001100110011000100010011000000;
LUT6 ii2170 (
	. xy ( \ii2170|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[6]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2170.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2170.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2170.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[0]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[0]|qx_net  ),
	. di ( \ii3344|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[10] .always_en = 1;
LUT6 ii2171 (
	. xy ( \ii2171|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[7]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2171.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2171.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2171.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1]|qx_net  ),
	. di ( \ii2595|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. di ( \ii2763|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[0] .always_en = 1;
LUT6 ii2172 (
	. xy ( \ii2172|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[8]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2172.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2172.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2172.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2173 (
	. xy ( \ii2173|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[9]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2173.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2173.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2173.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37]|qx_net  ),
	. di ( \ii2186|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .PLACE_LOCATION = "C18R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .PCK_LOCATION = "C18R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_10__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .PCK_LOCATION = "C18R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[4] .always_en = 1;
LUT6 ii2174 (
	. xy ( \ii2174|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[10]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2174.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2174.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2174.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .PLACE_LOCATION = "C10R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .PCK_LOCATION = "C10R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[3] .always_en = 1;
LUT6 ii2175 (
	. xy ( \ii2175|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[11]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2175.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2175.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2175.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
LUT6 ii2176 (
	. xy ( \ii2176|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[12]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2176.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.lut_0";
defparam ii2176.PCK_LOCATION = "C14R17.lp0.lut_0";
defparam ii2176.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]|qx_net  ),
	. di ( \ii2503|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .PLACE_LOCATION = "C14R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .PCK_LOCATION = "C14R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24] .always_en = 1;
LUT6 ii2177 (
	. xy ( \ii2177|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[13]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2177.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2177.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2177.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10]|qx_net  ),
	. di ( \ii2221|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10] .always_en = 0;
REG glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg|qx_net  ),
	. di ( \ii3312|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_hs_delay_en_reg.always_en = 1;
LUT6 ii2178 (
	. xy ( \ii2178|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2178.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2178.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2178.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2179 (
	. xy ( \ii2179|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[14]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2179.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2179.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2179.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2180 (
	. xy ( \ii2180|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[15]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2180.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2180.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2180.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[1]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[1]|qx_net  ),
	. di ( \ii3347|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[1] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[11] .always_en = 1;
LUT6 ii2181 (
	. xy ( \ii2181|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[16]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2181.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2181.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2181.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
ADD1_A carry_9_10__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_10__ADD_0|co_net  ),
	. s ( \carry_9_10__ADD_0|s_net  )
);
defparam carry_9_10__ADD_0.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_0.a_inv = "true";
defparam carry_9_10__ADD_0.PCK_LOCATION = "C18R11.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2]|qx_net  ),
	. di ( \ii2600|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .PLACE_LOCATION = "C18R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .PCK_LOCATION = "C18R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. di ( \ii2816|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[1] .always_en = 1;
LUT6 ii2182 (
	. xy ( \ii2182|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[17]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2182.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2182.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2182.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
ADD1_A carry_9_10__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[1]|qx_net  ),
	. ci ( \carry_9_10__ADD_0|co_net  ),
	. co ( \carry_9_10__ADD_1|co_net  ),
	. s ( \carry_9_10__ADD_1|s_net  )
);
defparam carry_9_10__ADD_1.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_1.a_inv = "true";
defparam carry_9_10__ADD_1.PCK_LOCATION = "C18R11.lp0.add2.add0";
LUT6 ii2183 (
	. xy ( \ii2183|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[18]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2183.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2183.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2183.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38]|qx_net  ),
	. di ( \ii2187|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38] .always_en = 0;
ADD1_A carry_9_10__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[2]|qx_net  ),
	. ci ( \carry_9_10__ADD_1|co_net  ),
	. co ( \carry_9_10__ADD_2|co_net  ),
	. s ( \carry_9_10__ADD_2|s_net  )
);
defparam carry_9_10__ADD_2.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_2.a_inv = "true";
defparam carry_9_10__ADD_2.PCK_LOCATION = "C18R11.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .PLACE_LOCATION = "C20R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .PCK_LOCATION = "C20R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_10__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[5] .always_en = 1;
LUT6 ii2184 (
	. xy ( \ii2184|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[19]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2184.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2184.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2184.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
ADD1_A carry_9_10__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[3]|qx_net  ),
	. ci ( \carry_9_10__ADD_2|co_net  ),
	. co ( \carry_9_10__ADD_3|co_net  ),
	. s ( \carry_9_10__ADD_3|s_net  )
);
defparam carry_9_10__ADD_3.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_3.a_inv = "true";
defparam carry_9_10__ADD_3.PCK_LOCATION = "C18R11.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .PLACE_LOCATION = "C14R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .PCK_LOCATION = "C14R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[4] .always_en = 1;
LUT6 ii2185 (
	. xy ( \ii2185|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[20]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2185.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2185.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2185.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
ADD1_A carry_9_10__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[4]|qx_net  ),
	. ci ( \carry_9_10__ADD_3|co_net  ),
	. co ( \carry_9_10__ADD_4|co_net  ),
	. s ( \carry_9_10__ADD_4|s_net  )
);
defparam carry_9_10__ADD_4.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_4.a_inv = "true";
defparam carry_9_10__ADD_4.PCK_LOCATION = "C18R11.lp0.add2.add0";
LUT6 ii2186 (
	. xy ( \ii2186|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2186.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2186.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2186.config_data = 64'b1111111111111111111111111111111111110000010100001111111101011100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]|qx_net  ),
	. di ( \ii2504|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[8] .always_en = 1;
ADD1_A carry_9_10__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[5]|qx_net  ),
	. ci ( \carry_9_10__ADD_4|co_net  ),
	. co ( \carry_9_10__ADD_5|co_net  ),
	. s ( \carry_9_10__ADD_5|s_net  )
);
defparam carry_9_10__ADD_5.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_5.a_inv = "true";
defparam carry_9_10__ADD_5.PCK_LOCATION = "C18R11.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25] .always_en = 1;
LUT6 ii2187 (
	. xy ( \ii2187|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[22]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2187.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2187.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2187.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11]|qx_net  ),
	. di ( \ii2222|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11] .always_en = 0;
ADD1_A carry_9_10__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[6]|qx_net  ),
	. ci ( \carry_9_10__ADD_5|co_net  ),
	. co ( \carry_9_10__ADD_6|co_net  ),
	. s ( \carry_9_10__ADD_6|s_net  )
);
defparam carry_9_10__ADD_6.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_6.a_inv = "true";
defparam carry_9_10__ADD_6.PCK_LOCATION = "C18R11.lp0.add2.add0";
LUT6 ii2188 (
	. xy ( \ii2188|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[23]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2188.PLACE_LOCATION = "C14R18.le_tile.le_guts.lp0.lut_0";
defparam ii2188.PCK_LOCATION = "C14R18.lp0.lut_0";
defparam ii2188.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
ADD1_A carry_9_10__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_9_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_8_reg[7]|qx_net  ),
	. ci ( \carry_9_10__ADD_6|co_net  ),
	. co ( \carry_9_10__ADD_7|co_net  ),
	. s ( \carry_9_10__ADD_7|s_net  )
);
defparam carry_9_10__ADD_7.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_7.a_inv = "true";
defparam carry_9_10__ADD_7.PCK_LOCATION = "C18R11.lp0.add2.add0";
LUT6 ii2189 (
	. xy ( \ii2189|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2189.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2189.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2189.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2190 (
	. xy ( \ii2190|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[24]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2190.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2190.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2190.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
LUT6 ii2200 (
	. xy ( \ii2200|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2200.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2200.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2200.config_data = 64'b0000000000000000101100111000000000000000000000001011001110000000;
REG mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg (
	. qx ( \mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg|qx_net  ),
	. di ( \ii3334|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.latch_mode = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.init = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.sr_inv = 1;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.sync_mode = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.no_sr = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.sr_value = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.PCK_LOCATION = "C4R16.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.clk_inv = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.en_inv = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HREADY_s_reg.always_en = 1;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[2]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[2]|qx_net  ),
	. di ( \ii3350|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[12] .always_en = 1;
ADD1_A carry_9_10__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_10__ADD_7|co_net  ),
	. co ( \carry_9_10__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_10__ADD_8.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_10__ADD_8.a_inv = "false";
defparam carry_9_10__ADD_8.PCK_LOCATION = "C18R12.lp0.add2.add0";
LUT6 ii2191 (
	. xy ( \ii2191|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[25]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2191.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2191.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2191.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
LUT6 ii2201 (
	. xy ( \ii2201|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[34]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2201.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2201.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2201.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3]|qx_net  ),
	. di ( \ii2601|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .PLACE_LOCATION = "C18R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .PCK_LOCATION = "C18R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. di ( \ii2849|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[2] .always_en = 1;
LUT6 ii2192 (
	. xy ( \ii2192|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[26]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2192.PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.lut_0";
defparam ii2192.PCK_LOCATION = "C14R20.lp0.lut_0";
defparam ii2192.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
LUT6 ii2202 (
	. xy ( \ii2202|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[35]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2202.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2202.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2202.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2193 (
	. xy ( \ii2193|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[27]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2193.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2193.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2193.config_data = 64'b0000000000000000000000000000000010101111000011111010001100000000;
LUT6 ii2203 (
	. xy ( \ii2203|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[36]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2203.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2203.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2203.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_reg_din_reg[0]  (
	. qx ( \mcu_arbiter_reg_din_reg[0]|qx_net  ),
	. di ( \ii3323|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[0] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[0] .init = 0;
defparam \mcu_arbiter_reg_din_reg[0] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[0] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[0] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[0] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[0] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[0] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[0] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[0] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[0] .always_en = 0;
LUT6 mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf.PLACE_LOCATION = "C10R13.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf.PCK_LOCATION = "C10R13.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40]|qx_net  ),
	. di ( \ii2190|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39]|qx_net  ),
	. di ( \ii2188|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .PCK_LOCATION = "C14R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_10__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[6] .always_en = 1;
LUT6 ii2194 (
	. xy ( \ii2194|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[28]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2194.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2194.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2194.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
LUT6 ii2204 (
	. xy ( \ii2204|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[37]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2204.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.lut_0";
defparam ii2204.PCK_LOCATION = "C14R22.lp0.lut_0";
defparam ii2204.config_data = 64'b0000110000001100000011000000110000000100000001000000110000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .PLACE_LOCATION = "C14R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .PCK_LOCATION = "C14R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[5] .always_en = 1;
LUT6 ii2195 (
	. xy ( \ii2195|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[29]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2195.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2195.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2195.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
LUT6 ii2205 (
	. xy ( \ii2205|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[38]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2205.PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.lut_0";
defparam ii2205.PCK_LOCATION = "C14R21.lp0.lut_0";
defparam ii2205.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2196 (
	. xy ( \ii2196|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[30]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2196.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2196.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2196.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
LUT6 ii2206 (
	. xy ( \ii2206|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[39]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2206.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2206.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2206.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[10]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[10]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[10] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]|qx_net  ),
	. di ( \ii2505|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .PCK_LOCATION = "C16R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .PLACE_LOCATION = "C16R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .PCK_LOCATION = "C16R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[0] .always_en = 1;
LUT6 ii2197 (
	. xy ( \ii2197|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[31]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2197.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.lut_0";
defparam ii2197.PCK_LOCATION = "C16R17.lp0.lut_0";
defparam ii2197.config_data = 64'b1111010011110100111101001111010011110100111101001111010011110100;
LUT6 ii2207 (
	. xy ( \ii2207|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[40]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2207.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2207.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2207.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12]|qx_net  ),
	. di ( \ii2223|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12] .always_en = 0;
REG glue_rd_start_s_reg (
	. qx ( \glue_rd_start_s_reg|qx_net  ),
	. di ( \glue_rd_start_f_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rd_start_s_reg.latch_mode = 0;
defparam glue_rd_start_s_reg.init = 0;
defparam glue_rd_start_s_reg.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam glue_rd_start_s_reg.sr_inv = 1;
defparam glue_rd_start_s_reg.sync_mode = 0;
defparam glue_rd_start_s_reg.no_sr = 0;
defparam glue_rd_start_s_reg.sr_value = 0;
defparam glue_rd_start_s_reg.PCK_LOCATION = "C16R17.lp0.reg0";
defparam glue_rd_start_s_reg.clk_inv = 0;
defparam glue_rd_start_s_reg.en_inv = 0;
defparam glue_rd_start_s_reg.always_en = 1;
LUT6 ii2198 (
	. xy ( \ii2198|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[32]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2198.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2198.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2198.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2208 (
	. xy ( \ii2208|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2208.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2208.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2208.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2199 (
	. xy ( \ii2199|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[33]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2199.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2199.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2199.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2209 (
	. xy ( \ii2209|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2209.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2209.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2209.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2210 (
	. xy ( \ii2210|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2210.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2210.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2210.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[3]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[3]|qx_net  ),
	. di ( \ii3353|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .PLACE_LOCATION = "C6R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .PCK_LOCATION = "C6R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[13] .always_en = 1;
LUT6 ii2211 (
	. xy ( \ii2211|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2211.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2211.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2211.config_data = 64'b0000000000000000000000000000000011111111010111111111110001011100;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4]|qx_net  ),
	. di ( \ii2602|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. di ( \ii2852|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[3] .always_en = 1;
LUT6 ii2212 (
	. xy ( \ii2212|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2212.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2212.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2212.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2213 (
	. xy ( \ii2213|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2213.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2213.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2213.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_reg_din_reg[1]  (
	. qx ( \mcu_arbiter_reg_din_reg[1]|qx_net  ),
	. di ( \ii3325|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[1] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[1] .init = 0;
defparam \mcu_arbiter_reg_din_reg[1] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[1] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[1] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[1] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[1] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[1] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[1] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[1] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[1] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41]|qx_net  ),
	. di ( \ii2191|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[41] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_10__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[7] .always_en = 1;
LUT6 ii2214 (
	. xy ( \ii2214|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2214.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2214.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2214.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .PLACE_LOCATION = "C10R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .PCK_LOCATION = "C10R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[6] .always_en = 1;
LUT6 ii2215 (
	. xy ( \ii2215|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2215.PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.lut_0";
defparam ii2215.PCK_LOCATION = "C16R18.lp0.lut_0";
defparam ii2215.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG glue_rx_packet_tx_packet_u_scaler_t9_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_sc1_fifo_readen_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.PCK_LOCATION = "C20R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t9_out1_reg.always_en = 1;
LUT6 ii2216 (
	. xy ( \ii2216|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2216.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2216.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2216.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[11]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[11]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[11] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]|qx_net  ),
	. di ( \ii2506|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0]|qx_net  ),
	. di ( \ii2381|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .PCK_LOCATION = "C8R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[1] .always_en = 1;
LUT6 ii2217 (
	. xy ( \ii2217|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2217.PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.lut_0";
defparam ii2217.PCK_LOCATION = "C16R22.lp0.lut_0";
defparam ii2217.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .PLACE_LOCATION = "C6R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .PCK_LOCATION = "C6R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13]|qx_net  ),
	. di ( \ii2224|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13] .always_en = 0;
LUT6 ii2218 (
	. xy ( \ii2218|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2218.PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.lut_0";
defparam ii2218.PCK_LOCATION = "C16R22.lp0.lut_0";
defparam ii2218.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2219 (
	. xy ( \ii2219|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2219.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2219.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2219.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2220 (
	. xy ( \ii2220|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2220.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.lut_0";
defparam ii2220.PCK_LOCATION = "C14R23.lp0.lut_0";
defparam ii2220.config_data = 64'b1100110011000000010001001100000011001100110000000100010011000000;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[4]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[4]|qx_net  ),
	. di ( \ii3356|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .PLACE_LOCATION = "C6R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .PCK_LOCATION = "C6R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[14] .always_en = 1;
LUT6 ii2221 (
	. xy ( \ii2221|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2221.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2221.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2221.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5]|qx_net  ),
	. di ( \ii2603|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. di ( \ii2855|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .PCK_LOCATION = "C14R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[4] .always_en = 1;
LUT6 ii2222 (
	. xy ( \ii2222|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2222.PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.lut_0";
defparam ii2222.PCK_LOCATION = "C16R22.lp0.lut_0";
defparam ii2222.config_data = 64'b1100110011001100010001001100000011001100110011000100010011000000;
LUT6 ii2223 (
	. xy ( \ii2223|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2223.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2223.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2223.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
REG \mcu_arbiter_reg_din_reg[2]  (
	. qx ( \mcu_arbiter_reg_din_reg[2]|qx_net  ),
	. di ( \ii3326|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[2] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[2] .init = 0;
defparam \mcu_arbiter_reg_din_reg[2] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[2] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[2] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[2] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[2] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[2] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[2] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[2] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42]|qx_net  ),
	. di ( \ii2192|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .PLACE_LOCATION = "C14R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .PCK_LOCATION = "C14R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[42] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8]|qx_net  ),
	. di ( \ii3253|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In2p_reg[8] .always_en = 1;
LUT6 ii2224 (
	. xy ( \ii2224|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[5]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2224.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2224.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2224.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .PLACE_LOCATION = "C14R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .PCK_LOCATION = "C14R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In3p_reg[7] .always_en = 1;
LUT6 ii2225 (
	. xy ( \ii2225|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[6]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2225.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2225.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2225.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2226 (
	. xy ( \ii2226|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[7]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2226.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2226.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2226.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[12]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[12]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[12] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]|qx_net  ),
	. di ( \ii2507|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1]|qx_net  ),
	. di ( \ii2411|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .PCK_LOCATION = "C8R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[2] .always_en = 1;
LUT6 ii2227 (
	. xy ( \ii2227|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[8]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2227.PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.lut_0";
defparam ii2227.PCK_LOCATION = "C16R22.lp0.lut_0";
defparam ii2227.config_data = 64'b1100110011001100010001001100000011001100110011000100010011000000;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .PLACE_LOCATION = "C6R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .PCK_LOCATION = "C6R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14]|qx_net  ),
	. di ( \ii2225|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .PCK_LOCATION = "C16R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14] .always_en = 0;
LUT6 ii2228 (
	. xy ( \ii2228|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[9]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2228.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2228.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2228.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
h6_r8051xc2 u_8051_u_h6_8051 (
	. clkcpu ( \u_pll_pll_u0|CO3_net  ),
	. clkper ( \u_pll_pll_u0|CO3_net  ),
	. hold ( \GND_0_inst|Y_net  ),
	. memack ( \ii2114|xy_net  ),
	. memdatai ( {
		/* memdatai [7] */ \ii2130|xy_net ,
		/* memdatai [6] */ \ii2128|xy_net ,
		/* memdatai [5] */ \ii2126|xy_net ,
		/* memdatai [4] */ \ii2124|xy_net ,
		/* memdatai [3] */ \ii2122|xy_net ,
		/* memdatai [2] */ \ii2120|xy_net ,
		/* memdatai [1] */ \ii2118|xy_net ,
		/* memdatai [0] */ \ii2116|xy_net 
	} ),
	. mempsack ( \ii2131|xy_net  ),
	. misoi ( ),
	. mosii ( ),
	. port0i ( {
		/* port0i [7] (nc) */ nc510 ,
		/* port0i [6] (nc) */ nc511 ,
		/* port0i [5] */ \io_phone_rst_inst|f_id[0]_net ,
		/* port0i [4] */ \ii2132|xy_net ,
		/* port0i [3] */ \glue_pasm_packet_finish_reg|qx_net ,
		/* port0i [2] (nc) */ nc512 ,
		/* port0i [1] (nc) */ nc513 ,
		/* port0i [0] (nc) */ nc514 
	} ),
	. port1i ( )
,
	. port2i ( )
,
	. port3i ( )
,
	. resetn ( \ii1982_dup|xy_net  ),
	. scki ( ),
	. scli ( ),
	. sdai ( ),
	. sfrack ( ),
	. sfrdatai ( )
,
	. ssn ( ),
	. swd ( ),
	. clkcpuen ( ),
	. clkperen ( ),
	. holda ( ),
	. intoccur ( ),
	. memaddr_comb ( {
		/* memaddr_comb [22] */ \u_8051_u_h6_8051|memaddr_comb[22]_net ,
		/* memaddr_comb [21] */ \u_8051_u_h6_8051|memaddr_comb[21]_net ,
		/* memaddr_comb [20] */ \u_8051_u_h6_8051|memaddr_comb[20]_net ,
		/* memaddr_comb [19] */ \u_8051_u_h6_8051|memaddr_comb[19]_net ,
		/* memaddr_comb [18] */ \u_8051_u_h6_8051|memaddr_comb[18]_net ,
		/* memaddr_comb [17] */ \u_8051_u_h6_8051|memaddr_comb[17]_net ,
		/* memaddr_comb [16] */ \u_8051_u_h6_8051|memaddr_comb[16]_net ,
		/* memaddr_comb [15] */ \u_8051_u_h6_8051|memaddr_comb[15]_net ,
		/* memaddr_comb [14] */ \u_8051_u_h6_8051|memaddr_comb[14]_net ,
		/* memaddr_comb [13] */ \u_8051_u_h6_8051|memaddr_comb[13]_net ,
		/* memaddr_comb [12] */ \u_8051_u_h6_8051|memaddr_comb[12]_net ,
		/* memaddr_comb [11] */ \u_8051_u_h6_8051|memaddr_comb[11]_net ,
		/* memaddr_comb [10] */ \u_8051_u_h6_8051|memaddr_comb[10]_net ,
		/* memaddr_comb [9] */ \u_8051_u_h6_8051|memaddr_comb[9]_net ,
		/* memaddr_comb [8] */ \u_8051_u_h6_8051|memaddr_comb[8]_net ,
		/* memaddr_comb [7] */ \u_8051_u_h6_8051|memaddr_comb[7]_net ,
		/* memaddr_comb [6] */ \u_8051_u_h6_8051|memaddr_comb[6]_net ,
		/* memaddr_comb [5] */ \u_8051_u_h6_8051|memaddr_comb[5]_net ,
		/* memaddr_comb [4] */ \u_8051_u_h6_8051|memaddr_comb[4]_net ,
		/* memaddr_comb [3] */ \u_8051_u_h6_8051|memaddr_comb[3]_net ,
		/* memaddr_comb [2] */ \u_8051_u_h6_8051|memaddr_comb[2]_net ,
		/* memaddr_comb [1] */ \u_8051_u_h6_8051|memaddr_comb[1]_net ,
		/* memaddr_comb [0] */ \u_8051_u_h6_8051|memaddr_comb[0]_net 
	} ),
	. memdatao_comb ( {
		/* memdatao_comb [7] */ \u_8051_u_h6_8051|memdatao_comb[7]_net ,
		/* memdatao_comb [6] */ \u_8051_u_h6_8051|memdatao_comb[6]_net ,
		/* memdatao_comb [5] */ \u_8051_u_h6_8051|memdatao_comb[5]_net ,
		/* memdatao_comb [4] */ \u_8051_u_h6_8051|memdatao_comb[4]_net ,
		/* memdatao_comb [3] */ \u_8051_u_h6_8051|memdatao_comb[3]_net ,
		/* memdatao_comb [2] */ \u_8051_u_h6_8051|memdatao_comb[2]_net ,
		/* memdatao_comb [1] */ \u_8051_u_h6_8051|memdatao_comb[1]_net ,
		/* memdatao_comb [0] */ \u_8051_u_h6_8051|memdatao_comb[0]_net 
	} ),
	. mempsrd_comb ( \u_8051_u_h6_8051|mempsrd_comb_net  ),
	. mempswr_comb ( \u_8051_u_h6_8051|mempswr_comb_net  ),
	. memrd_comb ( \u_8051_u_h6_8051|memrd_comb_net  ),
	. memwr_comb ( \u_8051_u_h6_8051|memwr_comb_net  ),
	. misoo ( ),
	. misotri ( ),
	. mosio ( ),
	. mositri ( ),
	. port0o ( {
		/* port0o [7] (nc) */ nc515 ,
		/* port0o [6] (nc) */ nc516 ,
		/* port0o [5] (nc) */ nc517 ,
		/* port0o [4] (nc) */ nc518 ,
		/* port0o [3] (nc) */ nc519 ,
		/* port0o [2] */ \u_8051_u_h6_8051|port0o[2]_net ,
		/* port0o [1] */ \u_8051_u_h6_8051|port0o[1]_net ,
		/* port0o [0] */ \u_8051_u_h6_8051|port0o[0]_net 
	} ),
	. port1o ( )
,
	. port2o ( )
,
	. port3o ( )
,
	. ro ( ),
	. scko ( ),
	. scktri ( ),
	. sclo ( ),
	. sdao ( ),
	. sfraddr ( )
,
	. sfrdatao ( )
,
	. sfroe ( ),
	. sfrwe ( ),
	. spssn ( )
,
	. waitstaten ( )
);
defparam u_8051_u_h6_8051.PLACE_LOCATION = "C23R28.h6_mcu_wrap.h6_mcu";
defparam u_8051_u_h6_8051.PCK_LOCATION = "NONE";
defparam u_8051_u_h6_8051.program_file = "../51_rx_pinf_tx_pinf_1080_reverse/Objects/mipi_rx_pinf_tx_pinf_1080.hex";
LUT6 ii2229 (
	. xy ( \ii2229|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[10]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2229.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2229.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2229.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2230 (
	. xy ( \ii2230|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[11]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2230.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2230.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2230.config_data = 64'b1111111011111110111111101111111011111110111111101111111011111110;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[5]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[5]|qx_net  ),
	. di ( \ii3359|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .PLACE_LOCATION = "C6R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .PCK_LOCATION = "C6R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .PLACE_LOCATION = "C6R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .PCK_LOCATION = "C6R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[15] .always_en = 1;
LUT6 ii2231 (
	. xy ( \ii2231|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2231.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.lut_0";
defparam ii2231.PCK_LOCATION = "C16R24.lp0.lut_0";
defparam ii2231.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6]|qx_net  ),
	. di ( \ii2604|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. di ( \ii2859|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .PCK_LOCATION = "C14R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[5] .always_en = 1;
LUT6 ii2232 (
	. xy ( \ii2232|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[12]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2232.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.lut_0";
defparam ii2232.PCK_LOCATION = "C16R24.lp0.lut_0";
defparam ii2232.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
LUT6 ii2233 (
	. xy ( \ii2233|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[13]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2233.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2233.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2233.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_reg_din_reg[3]  (
	. qx ( \mcu_arbiter_reg_din_reg[3]|qx_net  ),
	. di ( \ii3327|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[3] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[3] .init = 0;
defparam \mcu_arbiter_reg_din_reg[3] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[3] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[3] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[3] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[3] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[3] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[3] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[3] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43]|qx_net  ),
	. di ( \ii2193|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[43] .always_en = 0;
LUT6 ii2234 (
	. xy ( \ii2234|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[14]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2234.PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.lut_0";
defparam ii2234.PCK_LOCATION = "C16R19.lp0.lut_0";
defparam ii2234.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t43_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7] .always_en = 1;
LUT6 ii2235 (
	. xy ( \ii2235|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2235.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2235.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2235.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2236 (
	. xy ( \ii2236|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2236.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2236.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2236.config_data = 64'b1111111011111110111111101111111011111110111111101111111011111110;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[13]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[13]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[13] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]|qx_net  ),
	. di ( \ii2508|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2]|qx_net  ),
	. di ( \ii2412|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t104_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t5_out1_1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[3] .always_en = 1;
LUT6 ii2237 (
	. xy ( \ii2237|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2237.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2237.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2237.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .PLACE_LOCATION = "C8R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .PCK_LOCATION = "C8R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15]|qx_net  ),
	. di ( \ii2226|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .PCK_LOCATION = "C16R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[15] .always_en = 0;
LUT6 ii2238 (
	. xy ( \ii2238|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2238.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2238.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2238.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2239 (
	. xy ( \ii2239|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2239.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.lut_0";
defparam ii2239.PCK_LOCATION = "C16R24.lp0.lut_0";
defparam ii2239.config_data = 64'b0000110000001100000011000000110000000100000001000000110000000000;
LUT6 ii2240 (
	. xy ( \ii2240|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2240.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2240.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2240.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[6]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[6]|qx_net  ),
	. di ( \ii3362|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .PLACE_LOCATION = "C14R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .PCK_LOCATION = "C14R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[10] .always_en = 1;
LUT6 ii2241 (
	. xy ( \ii2241|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_fifo_empty_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2241.PLACE_LOCATION = "C16R25.le_tile.le_guts.lp0.lut_0";
defparam ii2241.PCK_LOCATION = "C16R25.lp0.lut_0";
defparam ii2241.config_data = 64'b0100010111001111010001011100111101000101110011110100010111001111;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7]|qx_net  ),
	. di ( \ii2605|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. di ( \ii2863|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[6] .always_en = 1;
LUT6 ii2242 (
	. xy ( \ii2242|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_hsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f0 ( \ii2241|xy_net  )
);
defparam ii2242.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2242.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2242.config_data = 64'b0000000000000000000000000000000001011111010111110101001101010000;
LUT6 ii2243 (
	. xy ( \ii2243|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2243.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.lut_0";
defparam ii2243.PCK_LOCATION = "C16R24.lp0.lut_0";
defparam ii2243.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \mcu_arbiter_reg_din_reg[4]  (
	. qx ( \mcu_arbiter_reg_din_reg[4]|qx_net  ),
	. di ( \ii3328|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[4] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[4] .init = 0;
defparam \mcu_arbiter_reg_din_reg[4] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[4] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[4] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[4] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[4] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[4] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[4] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[4] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44]|qx_net  ),
	. di ( \ii2194|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .PCK_LOCATION = "C16R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[44] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[0] .always_en = 1;
LUT6 ii2244 (
	. xy ( \ii2244|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2244.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2244.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2244.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2245 (
	. xy ( \ii2245|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23]|qx_net  ),
	. f0 ( \ii2160|xy_net  )
);
defparam ii2245.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2245.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2245.config_data = 64'b0000010000000100000001000000010000000100000001000000010000000100;
LUT6 ii2246 (
	. xy ( \ii2246|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2246.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2246.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2246.config_data = 64'b1100110011000000010001001100000011001100110000000100010011000000;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[14]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[14]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[14] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]|qx_net  ),
	. di ( \ii2509|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3]|qx_net  ),
	. di ( \ii2413|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[4] .always_en = 1;
LUT6 ii2247 (
	. xy ( \ii2247|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_fifo_empty_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2247.PLACE_LOCATION = "C16R25.le_tile.le_guts.lp0.lut_0";
defparam ii2247.PCK_LOCATION = "C16R25.lp0.lut_0";
defparam ii2247.config_data = 64'b0000000000000000000000000000000010111010000000000011000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16]|qx_net  ),
	. di ( \ii2227|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .PCK_LOCATION = "C16R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[16] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_2_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .PLACE_LOCATION = "C10R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .PCK_LOCATION = "C10R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_0_[3] .always_en = 1;
LUT6 ii2248 (
	. xy ( \ii2248|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2248.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.lut_0";
defparam ii2248.PCK_LOCATION = "C16R24.lp0.lut_0";
defparam ii2248.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2249 (
	. xy ( \ii2249|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2249.PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.lut_0";
defparam ii2249.PCK_LOCATION = "C16R22.lp0.lut_0";
defparam ii2249.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
LUT6 ii2250 (
	. xy ( \ii2250|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2250.PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.lut_0";
defparam ii2250.PCK_LOCATION = "C16R22.lp0.lut_0";
defparam ii2250.config_data = 64'b0000000010000000000000001000000000000000100000000000000010000000;
REG \mcu_arbiter_u_emif2apb_memdatai_reg[7]  (
	. qx ( \mcu_arbiter_u_emif2apb_memdatai_reg[7]|qx_net  ),
	. di ( \ii3365|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3339|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .init = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .PLACE_LOCATION = "C6R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .PCK_LOCATION = "C6R18.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_memdatai_reg[7] .always_en = 0;
LUT6 u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly (
	. xy ( \u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly|xy_net  )
);
defparam u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.lut_0";
defparam u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly.PCK_LOCATION = "NONE";
defparam u0_mipi1_clkdly_genblk1_0__u_mipi_clkdly.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[11] .always_en = 1;
LUT6 ii2251 (
	. xy ( \ii2251|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[0]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_last_line_flag_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2152|xy_net  ),
	. f0 ( \ii2150|xy_net  )
);
defparam ii2251.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2251.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2251.config_data = 64'b0000110000001100000011000000110000000100000001000000110000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8]|qx_net  ),
	. di ( \ii2606|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In3p_reg[7] .always_en = 1;
LUT6 ii2252 (
	. xy ( \ii2252|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \ii2167|xy_net  ),
	. f1 ( \ii2150|xy_net  ),
	. f0 ( \ii2166|xy_net  )
);
defparam ii2252.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.lut_0";
defparam ii2252.PCK_LOCATION = "C16R24.lp0.lut_0";
defparam ii2252.config_data = 64'b1010100010101010101000001010000010101000101010101010000010100000;
LUT6 ii2253 (
	. xy ( \ii2253|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0]|qx_net  )
);
defparam ii2253.PLACE_LOCATION = "C16R25.le_tile.le_guts.lp0.lut_0";
defparam ii2253.PCK_LOCATION = "C16R25.lp0.lut_0";
defparam ii2253.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
REG \mcu_arbiter_reg_din_reg[5]  (
	. qx ( \mcu_arbiter_reg_din_reg[5]|qx_net  ),
	. di ( \ii3329|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[5] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[5] .init = 0;
defparam \mcu_arbiter_reg_din_reg[5] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[5] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[5] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[5] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[5] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[5] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[5] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[5] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45]|qx_net  ),
	. di ( \ii2195|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .PCK_LOCATION = "C16R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[45] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[1] .always_en = 1;
LUT6 ii2254 (
	. xy ( \ii2254|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. f2 ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. f1 ( \ii2143|xy_net  ),
	. f0 ( \ii1984|xy_net  )
);
defparam ii2254.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.lut_0";
defparam ii2254.PCK_LOCATION = "C14R24.lp0.lut_0";
defparam ii2254.config_data = 64'b1111111111111111100000000000000011111111111111111000000000000000;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[15]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[15]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[15] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]|qx_net  ),
	. di ( \ii2510|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .PCK_LOCATION = "C18R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4]|qx_net  ),
	. di ( \ii2414|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17]|qx_net  ),
	. di ( \ii2228|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .PCK_LOCATION = "C16R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[17] .always_en = 0;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[9]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf.PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf.PCK_LOCATION = "C14R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_rstsf_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_rstsf_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rstrf_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[12] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[24]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .PLACE_LOCATION = "C18R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .PCK_LOCATION = "C18R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9]|qx_net  ),
	. di ( \ii2607|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0]|qx_net  ),
	. di ( \ii3285|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0] .always_en = 1;
REG \mcu_arbiter_reg_din_reg[6]  (
	. qx ( \mcu_arbiter_reg_din_reg[6]|qx_net  ),
	. di ( \ii3330|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[6] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[6] .init = 0;
defparam \mcu_arbiter_reg_din_reg[6] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[6] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[6] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[6] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[6] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[6] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[6] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[6] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46]|qx_net  ),
	. di ( \ii2196|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .PCK_LOCATION = "C16R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[46] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[2] .always_en = 1;
SPRAM_16Kx32 mcu_arbiter_u_psram_u_psram (
	. addr ( {
		/* addr [13] */ \GND_0_inst|Y_net ,
		/* addr [12] */ \u_8051_u_h6_8051|memaddr_comb[14]_net ,
		/* addr [11] */ \u_8051_u_h6_8051|memaddr_comb[13]_net ,
		/* addr [10] */ \u_8051_u_h6_8051|memaddr_comb[12]_net ,
		/* addr [9] */ \u_8051_u_h6_8051|memaddr_comb[11]_net ,
		/* addr [8] */ \u_8051_u_h6_8051|memaddr_comb[10]_net ,
		/* addr [7] */ \u_8051_u_h6_8051|memaddr_comb[9]_net ,
		/* addr [6] */ \u_8051_u_h6_8051|memaddr_comb[8]_net ,
		/* addr [5] */ \u_8051_u_h6_8051|memaddr_comb[7]_net ,
		/* addr [4] */ \u_8051_u_h6_8051|memaddr_comb[6]_net ,
		/* addr [3] */ \u_8051_u_h6_8051|memaddr_comb[5]_net ,
		/* addr [2] */ \u_8051_u_h6_8051|memaddr_comb[4]_net ,
		/* addr [1] */ \u_8051_u_h6_8051|memaddr_comb[3]_net ,
		/* addr [0] */ \u_8051_u_h6_8051|memaddr_comb[2]_net 
	} ),
	. beb ( {
		/* beb [3] */ \ii2044|xy_net ,
		/* beb [2] */ \ii2043|xy_net ,
		/* beb [1] */ \ii2042|xy_net ,
		/* beb [0] */ \ii2041|xy_net 
	} ),
	. ceb ( \ii2046|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  ),
	. datai ( {
		/* datai [31] */ \u_8051_u_h6_8051|memdatao_comb[7]_net ,
		/* datai [30] */ \u_8051_u_h6_8051|memdatao_comb[6]_net ,
		/* datai [29] */ \u_8051_u_h6_8051|memdatao_comb[5]_net ,
		/* datai [28] */ \u_8051_u_h6_8051|memdatao_comb[4]_net ,
		/* datai [27] */ \u_8051_u_h6_8051|memdatao_comb[3]_net ,
		/* datai [26] */ \u_8051_u_h6_8051|memdatao_comb[2]_net ,
		/* datai [25] */ \u_8051_u_h6_8051|memdatao_comb[1]_net ,
		/* datai [24] */ \u_8051_u_h6_8051|memdatao_comb[0]_net ,
		/* datai [23] */ \u_8051_u_h6_8051|memdatao_comb[7]_net ,
		/* datai [22] */ \u_8051_u_h6_8051|memdatao_comb[6]_net ,
		/* datai [21] */ \u_8051_u_h6_8051|memdatao_comb[5]_net ,
		/* datai [20] */ \u_8051_u_h6_8051|memdatao_comb[4]_net ,
		/* datai [19] */ \u_8051_u_h6_8051|memdatao_comb[3]_net ,
		/* datai [18] */ \u_8051_u_h6_8051|memdatao_comb[2]_net ,
		/* datai [17] */ \u_8051_u_h6_8051|memdatao_comb[1]_net ,
		/* datai [16] */ \u_8051_u_h6_8051|memdatao_comb[0]_net ,
		/* datai [15] */ \u_8051_u_h6_8051|memdatao_comb[7]_net ,
		/* datai [14] */ \u_8051_u_h6_8051|memdatao_comb[6]_net ,
		/* datai [13] */ \u_8051_u_h6_8051|memdatao_comb[5]_net ,
		/* datai [12] */ \u_8051_u_h6_8051|memdatao_comb[4]_net ,
		/* datai [11] */ \u_8051_u_h6_8051|memdatao_comb[3]_net ,
		/* datai [10] */ \u_8051_u_h6_8051|memdatao_comb[2]_net ,
		/* datai [9] */ \u_8051_u_h6_8051|memdatao_comb[1]_net ,
		/* datai [8] */ \u_8051_u_h6_8051|memdatao_comb[0]_net ,
		/* datai [7] */ \u_8051_u_h6_8051|memdatao_comb[7]_net ,
		/* datai [6] */ \u_8051_u_h6_8051|memdatao_comb[6]_net ,
		/* datai [5] */ \u_8051_u_h6_8051|memdatao_comb[5]_net ,
		/* datai [4] */ \u_8051_u_h6_8051|memdatao_comb[4]_net ,
		/* datai [3] */ \u_8051_u_h6_8051|memdatao_comb[3]_net ,
		/* datai [2] */ \u_8051_u_h6_8051|memdatao_comb[2]_net ,
		/* datai [1] */ \u_8051_u_h6_8051|memdatao_comb[1]_net ,
		/* datai [0] */ \u_8051_u_h6_8051|memdatao_comb[0]_net 
	} ),
	. web ( \ii2047|xy_net  ),
	. datao ( {
		/* datao [31] */ \mcu_arbiter_u_psram_u_psram|datao[31]_net ,
		/* datao [30] */ \mcu_arbiter_u_psram_u_psram|datao[30]_net ,
		/* datao [29] */ \mcu_arbiter_u_psram_u_psram|datao[29]_net ,
		/* datao [28] */ \mcu_arbiter_u_psram_u_psram|datao[28]_net ,
		/* datao [27] */ \mcu_arbiter_u_psram_u_psram|datao[27]_net ,
		/* datao [26] */ \mcu_arbiter_u_psram_u_psram|datao[26]_net ,
		/* datao [25] */ \mcu_arbiter_u_psram_u_psram|datao[25]_net ,
		/* datao [24] */ \mcu_arbiter_u_psram_u_psram|datao[24]_net ,
		/* datao [23] */ \mcu_arbiter_u_psram_u_psram|datao[23]_net ,
		/* datao [22] */ \mcu_arbiter_u_psram_u_psram|datao[22]_net ,
		/* datao [21] */ \mcu_arbiter_u_psram_u_psram|datao[21]_net ,
		/* datao [20] */ \mcu_arbiter_u_psram_u_psram|datao[20]_net ,
		/* datao [19] */ \mcu_arbiter_u_psram_u_psram|datao[19]_net ,
		/* datao [18] */ \mcu_arbiter_u_psram_u_psram|datao[18]_net ,
		/* datao [17] */ \mcu_arbiter_u_psram_u_psram|datao[17]_net ,
		/* datao [16] */ \mcu_arbiter_u_psram_u_psram|datao[16]_net ,
		/* datao [15] */ \mcu_arbiter_u_psram_u_psram|datao[15]_net ,
		/* datao [14] */ \mcu_arbiter_u_psram_u_psram|datao[14]_net ,
		/* datao [13] */ \mcu_arbiter_u_psram_u_psram|datao[13]_net ,
		/* datao [12] */ \mcu_arbiter_u_psram_u_psram|datao[12]_net ,
		/* datao [11] */ \mcu_arbiter_u_psram_u_psram|datao[11]_net ,
		/* datao [10] */ \mcu_arbiter_u_psram_u_psram|datao[10]_net ,
		/* datao [9] */ \mcu_arbiter_u_psram_u_psram|datao[9]_net ,
		/* datao [8] */ \mcu_arbiter_u_psram_u_psram|datao[8]_net ,
		/* datao [7] */ \mcu_arbiter_u_psram_u_psram|datao[7]_net ,
		/* datao [6] */ \mcu_arbiter_u_psram_u_psram|datao[6]_net ,
		/* datao [5] */ \mcu_arbiter_u_psram_u_psram|datao[5]_net ,
		/* datao [4] */ \mcu_arbiter_u_psram_u_psram|datao[4]_net ,
		/* datao [3] */ \mcu_arbiter_u_psram_u_psram|datao[3]_net ,
		/* datao [2] */ \mcu_arbiter_u_psram_u_psram|datao[2]_net ,
		/* datao [1] */ \mcu_arbiter_u_psram_u_psram|datao[1]_net ,
		/* datao [0] */ \mcu_arbiter_u_psram_u_psram|datao[0]_net 
	} )
);
defparam mcu_arbiter_u_psram_u_psram.PLACE_LOCATION = "C23R30.spram_16kx32_wrap.spram_16kx32";
defparam mcu_arbiter_u_psram_u_psram.PCK_LOCATION = "NONE";
defparam mcu_arbiter_u_psram_u_psram.init_file = "";
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[16]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[16]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .PLACE_LOCATION = "C4R15.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .PCK_LOCATION = "C4R15.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[16] .always_en = 0;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5]|qx_net  ),
	. di ( \ii2415|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18]|qx_net  ),
	. di ( \ii2229|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .PCK_LOCATION = "C16R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[18] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_rstsf_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_rstsf_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rstsf_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rstsf_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .PCK_LOCATION = "C16R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[13] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[25]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1]|qx_net  ),
	. di ( \ii3304|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1] .always_en = 1;
REG \mcu_arbiter_reg_din_reg[7]  (
	. qx ( \mcu_arbiter_reg_din_reg[7]|qx_net  ),
	. di ( \ii3331|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3324|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_reg_din_reg[7] .latch_mode = 0;
defparam \mcu_arbiter_reg_din_reg[7] .init = 0;
defparam \mcu_arbiter_reg_din_reg[7] .PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[7] .sr_inv = 1;
defparam \mcu_arbiter_reg_din_reg[7] .sync_mode = 0;
defparam \mcu_arbiter_reg_din_reg[7] .no_sr = 0;
defparam \mcu_arbiter_reg_din_reg[7] .sr_value = 0;
defparam \mcu_arbiter_reg_din_reg[7] .PCK_LOCATION = "C4R18.lp0.reg0";
defparam \mcu_arbiter_reg_din_reg[7] .clk_inv = 0;
defparam \mcu_arbiter_reg_din_reg[7] .en_inv = 0;
defparam \mcu_arbiter_reg_din_reg[7] .always_en = 0;
FIFO18K glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst (
	. dout ( {
		/* dout [63] (nc) */ nc520 ,
		/* dout [62] (nc) */ nc521 ,
		/* dout [61] (nc) */ nc522 ,
		/* dout [60] (nc) */ nc523 ,
		/* dout [59] (nc) */ nc524 ,
		/* dout [58] (nc) */ nc525 ,
		/* dout [57] (nc) */ nc526 ,
		/* dout [56] (nc) */ nc527 ,
		/* dout [55] (nc) */ nc528 ,
		/* dout [54] (nc) */ nc529 ,
		/* dout [53] (nc) */ nc530 ,
		/* dout [52] (nc) */ nc531 ,
		/* dout [51] (nc) */ nc532 ,
		/* dout [50] (nc) */ nc533 ,
		/* dout [49] (nc) */ nc534 ,
		/* dout [48] (nc) */ nc535 ,
		/* dout [47] (nc) */ nc536 ,
		/* dout [46] (nc) */ nc537 ,
		/* dout [45] (nc) */ nc538 ,
		/* dout [44] (nc) */ nc539 ,
		/* dout [43] (nc) */ nc540 ,
		/* dout [42] (nc) */ nc541 ,
		/* dout [41] (nc) */ nc542 ,
		/* dout [40] (nc) */ nc543 ,
		/* dout [39] (nc) */ nc544 ,
		/* dout [38] (nc) */ nc545 ,
		/* dout [37] (nc) */ nc546 ,
		/* dout [36] (nc) */ nc547 ,
		/* dout [35] (nc) */ nc548 ,
		/* dout [34] (nc) */ nc549 ,
		/* dout [33] (nc) */ nc550 ,
		/* dout [32] (nc) */ nc551 ,
		/* dout [31] (nc) */ nc552 ,
		/* dout [30] (nc) */ nc553 ,
		/* dout [29] (nc) */ nc554 ,
		/* dout [28] (nc) */ nc555 ,
		/* dout [27] (nc) */ nc556 ,
		/* dout [26] (nc) */ nc557 ,
		/* dout [25] (nc) */ nc558 ,
		/* dout [24] (nc) */ nc559 ,
		/* dout [23] (nc) */ nc560 ,
		/* dout [22] (nc) */ nc561 ,
		/* dout [21] (nc) */ nc562 ,
		/* dout [20] (nc) */ nc563 ,
		/* dout [19] (nc) */ nc564 ,
		/* dout [18] (nc) */ nc565 ,
		/* dout [17] (nc) */ nc566 ,
		/* dout [16] (nc) */ nc567 ,
		/* dout [15] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[15]_net ,
		/* dout [14] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[14]_net ,
		/* dout [13] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[13]_net ,
		/* dout [12] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[12]_net ,
		/* dout [11] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[11]_net ,
		/* dout [10] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[10]_net ,
		/* dout [9] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[9]_net ,
		/* dout [8] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[8]_net ,
		/* dout [7] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[7]_net ,
		/* dout [6] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[6]_net ,
		/* dout [5] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[5]_net ,
		/* dout [4] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[4]_net ,
		/* dout [3] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[3]_net ,
		/* dout [2] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[2]_net ,
		/* dout [1] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[1]_net ,
		/* dout [0] */ \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[0]_net 
	} ),
	. doutp ( )
,
	. din ( {
		/* din [63] */ \GND_0_inst|Y_net ,
		/* din [62] */ \GND_0_inst|Y_net ,
		/* din [61] */ \GND_0_inst|Y_net ,
		/* din [60] */ \GND_0_inst|Y_net ,
		/* din [59] */ \GND_0_inst|Y_net ,
		/* din [58] */ \GND_0_inst|Y_net ,
		/* din [57] */ \GND_0_inst|Y_net ,
		/* din [56] */ \GND_0_inst|Y_net ,
		/* din [55] */ \GND_0_inst|Y_net ,
		/* din [54] */ \GND_0_inst|Y_net ,
		/* din [53] */ \GND_0_inst|Y_net ,
		/* din [52] */ \GND_0_inst|Y_net ,
		/* din [51] */ \GND_0_inst|Y_net ,
		/* din [50] */ \GND_0_inst|Y_net ,
		/* din [49] */ \GND_0_inst|Y_net ,
		/* din [48] */ \GND_0_inst|Y_net ,
		/* din [47] */ \GND_0_inst|Y_net ,
		/* din [46] */ \GND_0_inst|Y_net ,
		/* din [45] */ \GND_0_inst|Y_net ,
		/* din [44] */ \GND_0_inst|Y_net ,
		/* din [43] */ \GND_0_inst|Y_net ,
		/* din [42] */ \GND_0_inst|Y_net ,
		/* din [41] */ \GND_0_inst|Y_net ,
		/* din [40] */ \GND_0_inst|Y_net ,
		/* din [39] */ \GND_0_inst|Y_net ,
		/* din [38] */ \GND_0_inst|Y_net ,
		/* din [37] */ \GND_0_inst|Y_net ,
		/* din [36] */ \GND_0_inst|Y_net ,
		/* din [35] */ \GND_0_inst|Y_net ,
		/* din [34] */ \GND_0_inst|Y_net ,
		/* din [33] */ \GND_0_inst|Y_net ,
		/* din [32] */ \GND_0_inst|Y_net ,
		/* din [31] */ \GND_0_inst|Y_net ,
		/* din [30] */ \GND_0_inst|Y_net ,
		/* din [29] */ \GND_0_inst|Y_net ,
		/* din [28] */ \GND_0_inst|Y_net ,
		/* din [27] */ \GND_0_inst|Y_net ,
		/* din [26] */ \GND_0_inst|Y_net ,
		/* din [25] */ \GND_0_inst|Y_net ,
		/* din [24] */ \GND_0_inst|Y_net ,
		/* din [23] */ \GND_0_inst|Y_net ,
		/* din [22] */ \GND_0_inst|Y_net ,
		/* din [21] */ \GND_0_inst|Y_net ,
		/* din [20] */ \GND_0_inst|Y_net ,
		/* din [19] */ \GND_0_inst|Y_net ,
		/* din [18] */ \GND_0_inst|Y_net ,
		/* din [17] */ \GND_0_inst|Y_net ,
		/* din [16] */ \GND_0_inst|Y_net ,
		/* din [15] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31]|qx_net ,
		/* din [14] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30]|qx_net ,
		/* din [13] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29]|qx_net ,
		/* din [12] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28]|qx_net ,
		/* din [11] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27]|qx_net ,
		/* din [10] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26]|qx_net ,
		/* din [9] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25]|qx_net ,
		/* din [8] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24]|qx_net ,
		/* din [7] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23]|qx_net ,
		/* din [6] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22]|qx_net ,
		/* din [5] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21]|qx_net ,
		/* din [4] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[20]|qx_net ,
		/* din [3] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[19]|qx_net ,
		/* din [2] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[18]|qx_net ,
		/* din [1] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[17]|qx_net ,
		/* din [0] */ \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[16]|qx_net 
	} ),
	. dinp ( {
		/* dinp [7] */ \GND_0_inst|Y_net ,
		/* dinp [6] */ \GND_0_inst|Y_net ,
		/* dinp [5] */ \GND_0_inst|Y_net ,
		/* dinp [4] */ \GND_0_inst|Y_net ,
		/* dinp [3] */ \GND_0_inst|Y_net ,
		/* dinp [2] */ \GND_0_inst|Y_net ,
		/* dinp [1] */ \GND_0_inst|Y_net ,
		/* dinp [0] */ \GND_0_inst|Y_net 
	} ),
	. writeclk ( \u_pll_pll_u0|CO0_net  ),
	. readclk ( \u_pll_pll_u0|CO0_net  ),
	. writeen ( \ii1990|xy_net  ),
	. readen ( \ii1989|xy_net  ),
	. reset ( \ii1987|xy_net  ),
	. regce ( \VCC_0_inst|Y_net  ),
	. writesave ( \GND_0_inst|Y_net  ),
	. writedrop ( \GND_0_inst|Y_net  ),
	. full ( ),
	. empty ( ),
	. almostfull ( ),
	. almostempty ( ),
	. overflow ( ),
	. underflow ( ),
	. eccoutdberr ( ),
	. eccoutsberr ( ),
	. eccreadaddr ( )
,
	. eccindberr ( \GND_0_inst|Y_net  ),
	. eccinsberr ( \GND_0_inst|Y_net  ),
	. writedropflag ( )
);
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.eccwriteen = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.writeclk_inv = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.eccreaden = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.readclk_inv = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.use_parity = 0;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.outreg = 1;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.almostfullth = 988;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.almostemptyth = 512;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.writewidth = 18;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.readwidth = 18;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.peek = 1;
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.PLACE_LOCATION = "C12R5.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
defparam glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst.PCK_LOCATION = "C12R5.u0_emb_top.emb18k_wrapper.u0_emb18k_core";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47]|qx_net  ),
	. di ( \ii2197|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .PCK_LOCATION = "C16R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[47] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[3] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[17]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[17]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[17] .always_en = 0;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6]|qx_net  ),
	. di ( \ii2416|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In3p_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20]|qx_net  ),
	. di ( \ii2232|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .PCK_LOCATION = "C16R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[20] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19]|qx_net  ),
	. di ( \ii2230|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .PCK_LOCATION = "C16R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[19] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[21] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[14] .always_en = 1;
LUT6 ii2281 (
	. xy ( \ii2281|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_10|s_net  )
);
defparam ii2281.PLACE_LOCATION = "C16R25.le_tile.le_guts.lp0.lut_0";
defparam ii2281.PCK_LOCATION = "C16R25.lp0.lut_0";
defparam ii2281.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[26]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_6__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2]|qx_net  ),
	. di ( \ii3305|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2] .always_en = 1;
LUT6 ii2282 (
	. xy ( \ii2282|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_11|s_net  )
);
defparam ii2282.PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.lut_0";
defparam ii2282.PCK_LOCATION = "C16R23.lp0.lut_0";
defparam ii2282.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[0] .always_en = 1;
REG glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg|qx_net  ),
	. di ( \ii3283|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_line_flag_reg.always_en = 1;
LUT6 ii2283 (
	. xy ( \ii2283|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_1|s_net  )
);
defparam ii2283.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2283.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2283.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48]|qx_net  ),
	. di ( \ii2198|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[48] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[4] .always_en = 1;
LUT6 ii2284 (
	. xy ( \ii2284|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_2|s_net  )
);
defparam ii2284.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2284.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2284.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[0]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2285 (
	. xy ( \ii2285|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_3|s_net  )
);
defparam ii2285.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2285.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2285.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2286 (
	. xy ( \ii2286|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_4|s_net  )
);
defparam ii2286.PLACE_LOCATION = "C16R20.le_tile.le_guts.lp0.lut_0";
defparam ii2286.PCK_LOCATION = "C16R20.lp0.lut_0";
defparam ii2286.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[18]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[18]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[10]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[18] .always_en = 0;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7]|qx_net  ),
	. di ( \ii2417|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .PCK_LOCATION = "C18R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7] .always_en = 0;
LUT6 ii2287 (
	. xy ( \ii2287|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_5|s_net  )
);
defparam ii2287.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2287.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2287.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21]|qx_net  ),
	. di ( \ii2233|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .PCK_LOCATION = "C16R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[21] .always_en = 0;
LUT6 ii2288 (
	. xy ( \ii2288|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_6|s_net  )
);
defparam ii2288.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2288.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2288.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2289 (
	. xy ( \ii2289|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_7|s_net  )
);
defparam ii2289.PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.lut_0";
defparam ii2289.PCK_LOCATION = "C16R21.lp0.lut_0";
defparam ii2289.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2290 (
	. xy ( \ii2290|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_8|s_net  )
);
defparam ii2290.PLACE_LOCATION = "C16R25.le_tile.le_guts.lp0.lut_0";
defparam ii2290.PCK_LOCATION = "C16R25.lp0.lut_0";
defparam ii2290.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2300 (
	. xy ( \ii2300|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8]|qx_net  ),
	. f0 ( \ii2299|xy_net  )
);
defparam ii2300.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.lut_0";
defparam ii2300.PCK_LOCATION = "C8R5.lp0.lut_0";
defparam ii2300.config_data = 64'b0100000001000000010000000100000001000000010000000100000001000000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[23]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[22] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[15] .always_en = 1;
LUT6 ii2291 (
	. xy ( \ii2291|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_sync_delay_vsync_dly_reg|qx_net  ),
	. f0 ( \carry_12_ADD_9|s_net  )
);
defparam ii2291.PLACE_LOCATION = "C16R25.le_tile.le_guts.lp0.lut_0";
defparam ii2291.PCK_LOCATION = "C16R25.lp0.lut_0";
defparam ii2291.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2301 (
	. xy ( \ii2301|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f1 ( \ii2300|xy_net  ),
	. f0 ( \ii2298|xy_net  )
);
defparam ii2301.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.lut_0";
defparam ii2301.PCK_LOCATION = "C10R5.lp0.lut_0";
defparam ii2301.config_data = 64'b1111000011110000111100001111101111110000111100001111000011110000;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[27]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .PCK_LOCATION = "C18R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_6__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3]|qx_net  ),
	. di ( \ii3306|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3] .always_en = 1;
LUT6 ii2292 (
	. xy ( \ii2292|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_flag_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_ack_d_reg|qx_net  ),
	. f1 ( \ii2167|xy_net  ),
	. f0 ( \ii2143|xy_net  )
);
defparam ii2292.PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.lut_0";
defparam ii2292.PCK_LOCATION = "C16R26.lp0.lut_0";
defparam ii2292.config_data = 64'b1101111111001100110111111100110011011111110011001101111111001100;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[1] .always_en = 1;
LUT6 ii2293 (
	. xy ( \ii2293|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_rx_cmd_valid_d_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_active_hs_d_reg|qx_net  )
);
defparam ii2293.PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.lut_0";
defparam ii2293.PCK_LOCATION = "C4R7.lp0.lut_0";
defparam ii2293.config_data = 64'b0000000000000000000000000000100000000000000000000000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50]|qx_net  ),
	. di ( \ii2201|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[50] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49]|qx_net  ),
	. di ( \ii2199|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .PCK_LOCATION = "C14R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[49] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_In1p_reg[5] .always_en = 1;
LUT6 ii2294 (
	. xy ( \ii2294|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[5]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[4]|qx_net  ),
	. f0 ( \ii2293|xy_net  )
);
defparam ii2294.PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.lut_0";
defparam ii2294.PCK_LOCATION = "C6R6.lp0.lut_0";
defparam ii2294.config_data = 64'b0010100000101000001010000010100000101000001010000010100000101000;
REG glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd_valid_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.PCK_LOCATION = "C4R8.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg.always_en = 1;
LUT6 ii2295 (
	. xy ( \ii2295|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[5]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_cmd_d_reg[4]|qx_net  ),
	. f0 ( \ii2293|xy_net  )
);
defparam ii2295.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.lut_0";
defparam ii2295.PCK_LOCATION = "C8R5.lp0.lut_0";
defparam ii2295.config_data = 64'b0000001000000010000000100000001000000010000000100000001000000010;
ADD1_A carry_9_7__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_7__ADD_0|co_net  ),
	. s ( \carry_9_7__ADD_0|s_net  )
);
defparam carry_9_7__ADD_0.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_0.a_inv = "true";
defparam carry_9_7__ADD_0.PCK_LOCATION = "C18R15.lp0.add2.add0";
LUT6 ii2296 (
	. xy ( \ii2296|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  )
);
defparam ii2296.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2296.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2296.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[19]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[19]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[11]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[19] .always_en = 0;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[20]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[20]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[12]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[20] .always_en = 0;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8]|qx_net  ),
	. di ( \ii2418|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8] .always_en = 0;
ADD1_A carry_9_7__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1]|qx_net  ),
	. ci ( \carry_9_7__ADD_0|co_net  ),
	. co ( \carry_9_7__ADD_1|co_net  ),
	. s ( \carry_9_7__ADD_1|s_net  )
);
defparam carry_9_7__ADD_1.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_1.a_inv = "true";
defparam carry_9_7__ADD_1.PCK_LOCATION = "C18R15.lp0.add2.add0";
LUT6 ii2297 (
	. xy ( \ii2297|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1]|qx_net  )
);
defparam ii2297.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2297.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2297.config_data = 64'b1111111111100000000000000000000011111111111000000000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22]|qx_net  ),
	. di ( \ii2234|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .PCK_LOCATION = "C16R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[22] .always_en = 0;
ADD1_A carry_9_7__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2]|qx_net  ),
	. ci ( \carry_9_7__ADD_1|co_net  ),
	. co ( \carry_9_7__ADD_2|co_net  ),
	. s ( \carry_9_7__ADD_2|s_net  )
);
defparam carry_9_7__ADD_2.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_2.a_inv = "true";
defparam carry_9_7__ADD_2.PCK_LOCATION = "C18R15.lp0.add2.add0";
LUT6 ii2298 (
	. xy ( \ii2298|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6]|qx_net  ),
	. f0 ( \ii2297|xy_net  )
);
defparam ii2298.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2298.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2298.config_data = 64'b0000000100000001000000010000000100000001000000010000000100000001;
ADD1_A carry_9_7__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3]|qx_net  ),
	. ci ( \carry_9_7__ADD_2|co_net  ),
	. co ( \carry_9_7__ADD_3|co_net  ),
	. s ( \carry_9_7__ADD_3|s_net  )
);
defparam carry_9_7__ADD_3.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_3.a_inv = "true";
defparam carry_9_7__ADD_3.PCK_LOCATION = "C18R15.lp0.add2.add0";
LUT6 ii2299 (
	. xy ( \ii2299|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0]|qx_net  )
);
defparam ii2299.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2299.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2299.config_data = 64'b0000000000000000000000000000000100000000000000000000000000000001;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[23] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4] .always_en = 1;
ADD1_A carry_9_7__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4]|qx_net  ),
	. ci ( \carry_9_7__ADD_3|co_net  ),
	. co ( \carry_9_7__ADD_4|co_net  ),
	. s ( \carry_9_7__ADD_4|s_net  )
);
defparam carry_9_7__ADD_4.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_4.a_inv = "true";
defparam carry_9_7__ADD_4.PCK_LOCATION = "C18R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .PLACE_LOCATION = "C4R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .PCK_LOCATION = "C4R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[16] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[28]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .PLACE_LOCATION = "C18R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .PCK_LOCATION = "C18R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4] .always_en = 1;
ADD1_A carry_9_7__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5]|qx_net  ),
	. ci ( \carry_9_7__ADD_4|co_net  ),
	. co ( \carry_9_7__ADD_5|co_net  ),
	. s ( \carry_9_7__ADD_5|s_net  )
);
defparam carry_9_7__ADD_5.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_5.a_inv = "true";
defparam carry_9_7__ADD_5.PCK_LOCATION = "C18R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_6__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4]|qx_net  ),
	. di ( \ii3307|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[2] .always_en = 1;
ADD1_A carry_9_7__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6]|qx_net  ),
	. ci ( \carry_9_7__ADD_5|co_net  ),
	. co ( \carry_9_7__ADD_6|co_net  ),
	. s ( \carry_9_7__ADD_6|s_net  )
);
defparam carry_9_7__ADD_6.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_6.a_inv = "true";
defparam carry_9_7__ADD_6.PCK_LOCATION = "C18R15.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51]|qx_net  ),
	. di ( \ii2202|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[51] .always_en = 0;
ADD1_A carry_9_7__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7]|qx_net  ),
	. ci ( \carry_9_7__ADD_6|co_net  ),
	. co ( \carry_9_7__ADD_7|co_net  ),
	. s ( \carry_9_7__ADD_7|s_net  )
);
defparam carry_9_7__ADD_7.PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_7.a_inv = "true";
defparam carry_9_7__ADD_7.PCK_LOCATION = "C18R15.lp0.add2.add0";
ADD1_A carry_9_7__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_7__ADD_7|co_net  ),
	. co ( \carry_9_7__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_7__ADD_8.PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_7__ADD_8.a_inv = "false";
defparam carry_9_7__ADD_8.PCK_LOCATION = "C18R16.lp0.add2.add0";
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[21]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[21]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[13]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[21] .always_en = 0;
REG \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9]|qx_net  ),
	. di ( \ii2419|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii1983|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .PCK_LOCATION = "C18R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .en_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23]|qx_net  ),
	. di ( \ii2235|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .PCK_LOCATION = "C16R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[23] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  ),
	. di ( \ii2578|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .PCK_LOCATION = "C8R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[24]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[24] .always_en = 1;
REG \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_cmd[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .PCK_LOCATION = "C10R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .PLACE_LOCATION = "C6R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .PCK_LOCATION = "C6R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[17] .always_en = 1;
REG glue_rx_packet_tx_packet_u_scaler_t86_out1_reg (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t86_out1_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.PLACE_LOCATION = "C6R20.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.sync_mode = 1;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.PCK_LOCATION = "C6R20.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_scaler_t86_out1_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[29]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_6__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5]|qx_net  ),
	. di ( \ii3308|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52]|qx_net  ),
	. di ( \ii2203|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[52] .always_en = 0;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[13]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[22]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[22]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[22] .always_en = 0;
PLLV2 u_pll_pll_u0 (
	. FBIN ( ),
	. FP_PLL_PDB ( ),
	. FP_PLL_RST ( ),
	. PLLCK0 ( \u_osc|OSC_net  ),
	. PLLCK1 ( ),
	. PSCK ( ),
	. PSDIR ( ),
	. PSEN ( ),
	. PSSEL ( )
,
	. fp_cf_clk ( ),
	. fp_cf_en ( ),
	. fp_cf_in ( ),
	. fp_cf_up ( ),
	. fp_cfg_sel ( ),
	. ACTIVECK ( ),
	. CKBAD0 ( ),
	. CKBAD1 ( ),
	. CO0 ( \u_pll_pll_u0|CO0_net  ),
	. CO1 ( \u_pll_pll_u0|CO1_net  ),
	. CO2 ( \u_pll_pll_u0|CO2_net  ),
	. CO3 ( \u_pll_pll_u0|CO3_net  ),
	. CO4 ( ),
	. CO5 ( ),
	. DTEST ( )
,
	. FBOUT ( ),
	. PLOCK ( \u_pll_pll_u0|PLOCK_net  ),
	. PSDONE ( ),
	. fp_cf_out ( )
);
defparam u_pll_pll_u0.CFG_DIVN = 7;
defparam u_pll_pll_u0.CFG_CO0DLY = 0;
defparam u_pll_pll_u0.CFG_FRAC = 2;
defparam u_pll_pll_u0.CFG_DTEST_EN = 0;
defparam u_pll_pll_u0.CFG_FP_EN = 0;
defparam u_pll_pll_u0.CFG_P4SEL = 2;
defparam u_pll_pll_u0.CFG_SSEN = 0;
defparam u_pll_pll_u0.CFG_BPS0 = 0;
defparam u_pll_pll_u0.CFG_CO3DLY = 0;
defparam u_pll_pll_u0.CFG_BPS1 = 0;
defparam u_pll_pll_u0.CFG_DIVC0 = 6;
defparam u_pll_pll_u0.PCK_LOCATION = "C24R25.pll";
defparam u_pll_pll_u0.CFG_DIVC1 = 74;
defparam u_pll_pll_u0.CFG_BPS2 = 0;
defparam u_pll_pll_u0.CFG_DIVC2 = 18;
defparam u_pll_pll_u0.CFG_BPS3 = 0;
defparam u_pll_pll_u0.CFG_DIVC3 = 24;
defparam u_pll_pll_u0.CFG_BPS4 = 0;
defparam u_pll_pll_u0.CFG_DIVC4 = 7;
defparam u_pll_pll_u0.CFG_RST_REG_ENB = 0;
defparam u_pll_pll_u0.CFG_BPS5 = 0;
defparam u_pll_pll_u0.CFG_DIVC5 = 8;
defparam u_pll_pll_u0.CFG_BP_VDOUT = 0;
defparam u_pll_pll_u0.CFG_ATEST_SEL = 0;
defparam u_pll_pll_u0.CFG_P2SEL = 0;
defparam u_pll_pll_u0.CFG_CP_AUTO_ENB = 0;
defparam u_pll_pll_u0.CFG_DTEST_SEL = 0;
defparam u_pll_pll_u0.CFG_PPDB_SEL = 1;
defparam u_pll_pll_u0.CFG_CALIB_RSTN = 1;
defparam u_pll_pll_u0.CFG_LKD_TOL = 0;
defparam u_pll_pll_u0.CFG_LPF = 2;
defparam u_pll_pll_u0.CFG_CKSEL = 0;
defparam u_pll_pll_u0.CFG_ATEST_EN = 0;
defparam u_pll_pll_u0.CFG_CO1DLY = 0;
defparam u_pll_pll_u0.CFG_BK = 1;
defparam u_pll_pll_u0.CFG_SEL_FBPATH = 0;
defparam u_pll_pll_u0.CFG_P5SEL = 0;
defparam u_pll_pll_u0.CFG_CK_SWITCH_EN = 0;
defparam u_pll_pll_u0.CFG_VCO_INI_SEL = 0;
defparam u_pll_pll_u0.CFG_CPSEL_CR = 2;
defparam u_pll_pll_u0.CFG_PFBSEL = 0;
defparam u_pll_pll_u0.CFG_P0SEL = 0;
defparam u_pll_pll_u0.CFG_LKD_MUX = 0;
defparam u_pll_pll_u0.CFG_CO4DLY = 6;
defparam u_pll_pll_u0.CFG_SSDIVH = 0;
defparam u_pll_pll_u0.CFG_MKEN0 = 1;
defparam u_pll_pll_u0.CFG_MKEN1 = 1;
defparam u_pll_pll_u0.CFG_SSDIVL = 99;
defparam u_pll_pll_u0.CFG_MKEN2 = 1;
defparam u_pll_pll_u0.CFG_MKEN3 = 1;
defparam u_pll_pll_u0.CFG_P3SEL = 0;
defparam u_pll_pll_u0.CFG_MKEN4 = 1;
defparam u_pll_pll_u0.CFG_CALIB_MANUAL = 8;
defparam u_pll_pll_u0.CFG_CALIB_WIN = 0;
defparam u_pll_pll_u0.CFG_MKEN5 = 0;
defparam u_pll_pll_u0.CFG_LKD_HOLD = 0;
defparam u_pll_pll_u0.CFG_CALIB_16_32U = 0;
defparam u_pll_pll_u0.CFG_RSTPLL_SEL = 1;
defparam u_pll_pll_u0.CFG_CO2DLY = 0;
defparam u_pll_pll_u0.CFG_CALIB_DIV = 10;
defparam u_pll_pll_u0.CFG_FORCE_LOCK = 0;
defparam u_pll_pll_u0.CFG_SSRG = 1;
defparam u_pll_pll_u0.CFG_LOCK_GATE = 1;
defparam u_pll_pll_u0.CFG_CPSEL_FN = 112;
defparam u_pll_pll_u0.CFG_FLDD = 3;
defparam u_pll_pll_u0.CFG_DIVFB = 0;
defparam u_pll_pll_u0.CFG_VRSEL = 2;
defparam u_pll_pll_u0.CFG_P1SEL = 0;
defparam u_pll_pll_u0.CFG_CALIB_EN = 1;
defparam u_pll_pll_u0.PLACE_LOCATION = "C24R25.array.C12R25.gclk_tile.c1r1_gclk_gen.pll";
defparam u_pll_pll_u0.CFG_CO5DLY = 0;
defparam u_pll_pll_u0.CFG_DIVM = 112;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24]|qx_net  ),
	. di ( \ii2236|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[24] .always_en = 0;
LUT6 ii2328 (
	. xy ( \ii2328|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_10|s_net  )
);
defparam ii2328.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.lut_0";
defparam ii2328.PCK_LOCATION = "C10R5.lp0.lut_0";
defparam ii2328.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. di ( \ii2580|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .PCK_LOCATION = "C8R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[0] .always_en = 1;
LUT6 ii2329 (
	. xy ( \ii2329|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_11|s_net  )
);
defparam ii2329.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.lut_0";
defparam ii2329.PCK_LOCATION = "C10R5.lp0.lut_0";
defparam ii2329.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2330 (
	. xy ( \ii2330|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_1|s_net  )
);
defparam ii2330.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2330.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2330.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[25]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[25] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .PLACE_LOCATION = "C8R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .PCK_LOCATION = "C8R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[18] .always_en = 1;
LUT6 ii2331 (
	. xy ( \ii2331|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_2|s_net  )
);
defparam ii2331.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2331.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2331.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[30]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_6__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6]|qx_net  ),
	. di ( \ii3309|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6] .always_en = 1;
LUT6 ii2332 (
	. xy ( \ii2332|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_3|s_net  )
);
defparam ii2332.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2332.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2332.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .PLACE_LOCATION = "C18R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .PCK_LOCATION = "C18R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0] .always_en = 1;
LUT6 ii2333 (
	. xy ( \ii2333|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_4|s_net  )
);
defparam ii2333.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2333.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2333.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53]|qx_net  ),
	. di ( \ii2204|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .PCK_LOCATION = "C16R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[53] .always_en = 0;
LUT6 ii2334 (
	. xy ( \ii2334|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_5|s_net  )
);
defparam ii2334.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2334.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2334.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2335 (
	. xy ( \ii2335|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_6|s_net  )
);
defparam ii2335.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2335.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2335.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2336 (
	. xy ( \ii2336|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_7|s_net  )
);
defparam ii2336.PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.lut_0";
defparam ii2336.PCK_LOCATION = "C8R4.lp0.lut_0";
defparam ii2336.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[23]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[23]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[23] .always_en = 0;
LUT6 ii2337 (
	. xy ( \ii2337|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_8|s_net  )
);
defparam ii2337.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.lut_0";
defparam ii2337.PCK_LOCATION = "C10R5.lp0.lut_0";
defparam ii2337.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25]|qx_net  ),
	. di ( \ii2237|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[25] .always_en = 0;
LUT6 ii2338 (
	. xy ( \ii2338|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  ),
	. f0 ( \carry_12_0__ADD_9|s_net  )
);
defparam ii2338.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.lut_0";
defparam ii2338.PCK_LOCATION = "C10R5.lp0.lut_0";
defparam ii2338.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. di ( \ii2583|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .PLACE_LOCATION = "C8R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .PCK_LOCATION = "C8R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[1] .always_en = 1;
LUT6 ii2339 (
	. xy ( \ii2339|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_sc1_rd_line_data_en_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10]|qx_net  ),
	. f0 ( \ii2298|xy_net  )
);
defparam ii2339.PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.lut_0";
defparam ii2339.PCK_LOCATION = "C10R5.lp0.lut_0";
defparam ii2339.config_data = 64'b0000001000000011000000110000001100000000000000000000000000000000;
LUT6 ii2340 (
	. xy ( \ii2340|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  )
);
defparam ii2340.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2340.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2340.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[26]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[26] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[20] .always_en = 1;
LUT6 ii2341 (
	. xy ( \ii2341|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_data_process_frame_start_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  )
);
defparam ii2341.PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.lut_0";
defparam ii2341.PCK_LOCATION = "C16R6.lp0.lut_0";
defparam ii2341.config_data = 64'b1110110011101100111011001110110011101100111011001110110011101100;
REG \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[31]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_6__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7]|qx_net  ),
	. di ( \ii3310|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_0_[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .PCK_LOCATION = "C8R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_1_[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54]|qx_net  ),
	. di ( \ii2205|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .PCK_LOCATION = "C16R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[54] .always_en = 0;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[24]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[24]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .PCK_LOCATION = "C6R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[24] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0]|qx_net  ),
	. di ( \ii2495|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .PCK_LOCATION = "C16R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26]|qx_net  ),
	. di ( \ii2238|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[26] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .PCK_LOCATION = "C16R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[27]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[27] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[21] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_6__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2] .always_en = 1;
REG mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg (
	. qx ( \mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg|qx_net  ),
	. di ( \ii3338|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.latch_mode = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.init = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.PLACE_LOCATION = "C6R14.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.sr_inv = 1;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.sync_mode = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.no_sr = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.sr_value = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.PCK_LOCATION = "C6R14.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.clk_inv = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.en_inv = 0;
defparam mcu_arbiter_u_emif2apb_fpga_HWRITE_reg_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55]|qx_net  ),
	. di ( \ii2206|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .PLACE_LOCATION = "C16R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .PCK_LOCATION = "C16R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[55] .always_en = 0;
ADD1_A carry_12_1__ADD_10 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10]|qx_net  ),
	. ci ( \carry_12_1__ADD_9|co_net  ),
	. co ( \carry_12_1__ADD_10|co_net  ),
	. s ( \carry_12_1__ADD_10|s_net  )
);
defparam carry_12_1__ADD_10.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_10.a_inv = "false";
defparam carry_12_1__ADD_10.PCK_LOCATION = "C18R5.lp0.add2.add0";
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[25]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[25]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[25] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[0]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[0]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1]|qx_net  ),
	. di ( \ii2496|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .PCK_LOCATION = "C16R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[1] .always_en = 1;
ADD1_A carry_12_1__ADD_11 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11]|qx_net  ),
	. ci ( \carry_12_1__ADD_10|co_net  ),
	. co ( ),
	. s ( \carry_12_1__ADD_11|s_net  )
);
defparam carry_12_1__ADD_11.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_1__ADD_11.a_inv = "false";
defparam carry_12_1__ADD_11.PCK_LOCATION = "C18R5.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27]|qx_net  ),
	. di ( \ii2239|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .PCK_LOCATION = "C14R25.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[27] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .PLACE_LOCATION = "C16R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .PCK_LOCATION = "C16R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[28]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[28] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[22] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_6__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56]|qx_net  ),
	. di ( \ii2207|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .PCK_LOCATION = "C16R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[56] .always_en = 0;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg|qx_net  ),
	. di ( \ii2145|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.PLACE_LOCATION = "C14R30.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.PCK_LOCATION = "C14R30.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_fifo_readen_generator_inst_is_3Eh_request_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[0] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[26]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[26]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[26] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[1]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[1]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2]|qx_net  ),
	. di ( \ii2497|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .PCK_LOCATION = "C16R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28]|qx_net  ),
	. di ( \ii2240|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[28] .always_en = 0;
LUT6 ii2368 (
	. xy ( \ii2368|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_10|s_net  )
);
defparam ii2368.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2368.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2368.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[4] .always_en = 1;
LUT6 ii2369 (
	. xy ( \ii2369|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_11|s_net  )
);
defparam ii2369.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2369.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2369.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2370 (
	. xy ( \ii2370|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_1|s_net  )
);
defparam ii2370.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2370.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2370.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0]|qx_net  ),
	. di ( \ii2556|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[30]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[30] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[29]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .PCK_LOCATION = "C8R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[23] .always_en = 1;
LUT6 ii2371 (
	. xy ( \ii2371|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_2|s_net  )
);
defparam ii2371.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2371.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2371.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8]|qx_net  ),
	. di ( \ii3137|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In2p_reg[8] .always_en = 1;
LUT6 ii2372 (
	. xy ( \ii2372|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_3|s_net  )
);
defparam ii2372.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2372.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2372.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4] .always_en = 1;
LUT6 ii2373 (
	. xy ( \ii2373|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_4|s_net  )
);
defparam ii2373.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2373.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2373.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57]|qx_net  ),
	. di ( \ii2208|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .PCK_LOCATION = "C14R23.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[57] .always_en = 0;
LUT6 ii2374 (
	. xy ( \ii2374|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_5|s_net  )
);
defparam ii2374.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2374.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2374.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2375 (
	. xy ( \ii2375|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_6|s_net  )
);
defparam ii2375.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2375.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2375.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[1] .always_en = 1;
LUT6 ii2376 (
	. xy ( \ii2376|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_7|s_net  )
);
defparam ii2376.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2376.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2376.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[27]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[27]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .PLACE_LOCATION = "C4R14.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .PCK_LOCATION = "C4R14.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[27] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[2]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[2]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3]|qx_net  ),
	. di ( \ii2498|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .PLACE_LOCATION = "C16R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .PCK_LOCATION = "C16R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_12__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[0] .always_en = 1;
LUT6 ii2377 (
	. xy ( \ii2377|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_8|s_net  )
);
defparam ii2377.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2377.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2377.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .PLACE_LOCATION = "C10R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .PCK_LOCATION = "C10R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30]|qx_net  ),
	. di ( \ii2244|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .PCK_LOCATION = "C16R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[30] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29]|qx_net  ),
	. di ( \ii2242|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .PCK_LOCATION = "C14R24.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[29] .always_en = 0;
LUT6 ii2378 (
	. xy ( \ii2378|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_2__ADD_9|s_net  )
);
defparam ii2378.PLACE_LOCATION = "C16R4.le_tile.le_guts.lp0.lut_0";
defparam ii2378.PCK_LOCATION = "C16R4.lp0.lut_0";
defparam ii2378.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[5] .always_en = 1;
LUT6 ii2379 (
	. xy ( \ii2379|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[8]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[7]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[6]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[5]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[4]|qx_net  )
);
defparam ii2379.PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.lut_0";
defparam ii2379.PCK_LOCATION = "C16R5.lp0.lut_0";
defparam ii2379.config_data = 64'b0000000000000000000000000000000000000000000000000000000001111111;
LUT6 ii2380 (
	. xy ( \ii2380|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_data_process_frame_start_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[11]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_rd_line_cnt_reg[10]|qx_net  ),
	. f0 ( \ii2379|xy_net  )
);
defparam ii2380.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2380.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2380.config_data = 64'b0010111100000000001011110000000000101111000000000010111100000000;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1]|qx_net  ),
	. di ( \ii2559|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_rx_payload_d_reg[31]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .PCK_LOCATION = "C8R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_data_process_fifo_din_reg[31] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[24]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[24] .always_en = 1;
LUT6 ii2381 (
	. xy ( \ii2381|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  )
);
defparam ii2381.PLACE_LOCATION = "C18R4.le_tile.le_guts.lp0.lut_0";
defparam ii2381.PCK_LOCATION = "C18R4.lp0.lut_0";
defparam ii2381.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58]|qx_net  ),
	. di ( \ii2209|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[58] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .PCK_LOCATION = "C8R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .PCK_LOCATION = "C18R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[2] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[28]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[28]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .PCK_LOCATION = "C4R13.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[28] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[3]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[3]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .PLACE_LOCATION = "C4R5.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .PCK_LOCATION = "C4R5.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4]|qx_net  ),
	. di ( \ii2499|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .PCK_LOCATION = "C18R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_12__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31]|qx_net  ),
	. di ( \ii2245|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .PCK_LOCATION = "C16R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_reg[31] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2]|qx_net  ),
	. di ( \ii2560|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[25]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[25] .always_en = 1;
REG mcu_arbiter_u_emif2apb_memrd_s_reg (
	. qx ( \mcu_arbiter_u_emif2apb_memrd_s_reg|qx_net  ),
	. di ( \ii3333|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.latch_mode = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.init = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.sr_inv = 1;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.sync_mode = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.no_sr = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.sr_value = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.PCK_LOCATION = "C4R16.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.clk_inv = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.en_inv = 0;
defparam mcu_arbiter_u_emif2apb_memrd_s_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0]|qx_net  ),
	. di ( \ii2430|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60]|qx_net  ),
	. di ( \ii2212|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .PLACE_LOCATION = "C14R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .PCK_LOCATION = "C14R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[60] .always_en = 0;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59]|qx_net  ),
	. di ( \ii2210|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .PLACE_LOCATION = "C16R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .PCK_LOCATION = "C16R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[59] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[3] .always_en = 1;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[29]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[29]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[21]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .PCK_LOCATION = "C4R13.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[29] .always_en = 0;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[30]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[30]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[22]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .PCK_LOCATION = "C4R13.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[30] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[4]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[4]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5]|qx_net  ),
	. di ( \ii2500|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .PCK_LOCATION = "C18R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_12__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In3p_reg[7] .always_en = 1;
LUT6 ii2409 (
	. xy ( \ii2409|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_10|s_net  )
);
defparam ii2409.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.lut_0";
defparam ii2409.PCK_LOCATION = "C18R5.lp0.lut_0";
defparam ii2409.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2410 (
	. xy ( \ii2410|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_11|s_net  )
);
defparam ii2410.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.lut_0";
defparam ii2410.PCK_LOCATION = "C18R5.lp0.lut_0";
defparam ii2410.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3]|qx_net  ),
	. di ( \ii2561|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[26]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[26] .always_en = 1;
LUT6 ii2411 (
	. xy ( \ii2411|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_1|s_net  )
);
defparam ii2411.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2411.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2411.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2412 (
	. xy ( \ii2412|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_2|s_net  )
);
defparam ii2412.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2412.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2412.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .PLACE_LOCATION = "C10R29.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .PCK_LOCATION = "C10R29.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7] .always_en = 1;
LUT6 ii2413 (
	. xy ( \ii2413|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_3|s_net  )
);
defparam ii2413.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2413.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2413.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61]|qx_net  ),
	. di ( \ii2213|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .PCK_LOCATION = "C16R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[61] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_11__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[0] .always_en = 1;
LUT6 ii2414 (
	. xy ( \ii2414|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_4|s_net  )
);
defparam ii2414.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2414.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2414.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2415 (
	. xy ( \ii2415|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_5|s_net  )
);
defparam ii2415.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2415.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2415.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .PCK_LOCATION = "C20R13.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[4] .always_en = 1;
LUT6 ii2416 (
	. xy ( \ii2416|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_6|s_net  )
);
defparam ii2416.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2416.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2416.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[5]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \mcu_arbiter_u_emif2apb_write_data_temp_reg[31]  (
	. qx ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[31]|qx_net  ),
	. di ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[23]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii3336|xy_net  ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .latch_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .init = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .PLACE_LOCATION = "C4R13.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .sr_inv = 1;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .sync_mode = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .no_sr = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .sr_value = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .PCK_LOCATION = "C4R13.lp0.reg0";
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .clk_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .en_inv = 0;
defparam \mcu_arbiter_u_emif2apb_write_data_temp_reg[31] .always_en = 0;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[5]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6]|qx_net  ),
	. di ( \ii2501|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10]|qx_net  ),
	. di ( \ii2328|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .PCK_LOCATION = "C10R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10] .always_en = 0;
ADD1_A carry_9_ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_ADD_0|co_net  ),
	. s ( \carry_9_ADD_0|s_net  )
);
defparam carry_9_ADD_0.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_0.a_inv = "true";
defparam carry_9_ADD_0.PCK_LOCATION = "C16R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_12__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[3] .always_en = 1;
LUT6 ii2417 (
	. xy ( \ii2417|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_7|s_net  )
);
defparam ii2417.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2417.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2417.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[3] .always_en = 1;
ADD1_A carry_9_ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[1]|qx_net  ),
	. ci ( \carry_9_ADD_0|co_net  ),
	. co ( \carry_9_ADD_1|co_net  ),
	. s ( \carry_9_ADD_1|s_net  )
);
defparam carry_9_ADD_1.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_1.a_inv = "true";
defparam carry_9_ADD_1.PCK_LOCATION = "C16R7.lp0.add2.add0";
LUT6 ii2418 (
	. xy ( \ii2418|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_8|s_net  )
);
defparam ii2418.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.lut_0";
defparam ii2418.PCK_LOCATION = "C18R5.lp0.lut_0";
defparam ii2418.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
ADD1_A carry_9_ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[2]|qx_net  ),
	. ci ( \carry_9_ADD_1|co_net  ),
	. co ( \carry_9_ADD_2|co_net  ),
	. s ( \carry_9_ADD_2|s_net  )
);
defparam carry_9_ADD_2.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_2.a_inv = "true";
defparam carry_9_ADD_2.PCK_LOCATION = "C16R7.lp0.add2.add0";
LUT6 ii2419 (
	. xy ( \ii2419|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \carry_12_1__ADD_9|s_net  )
);
defparam ii2419.PLACE_LOCATION = "C18R5.le_tile.le_guts.lp0.lut_0";
defparam ii2419.PCK_LOCATION = "C18R5.lp0.lut_0";
defparam ii2419.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2420 (
	. xy ( \ii2420|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[9]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[8]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[7]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[6]|qx_net  )
);
defparam ii2420.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2420.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2420.config_data = 64'b0000000000000001000000000000000100000000000000010000000000000001;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4]|qx_net  ),
	. di ( \ii2562|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4] .always_en = 1;
ADD1_A carry_13_ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_13_ADD_0|co_net  ),
	. s ( )
);
defparam carry_13_ADD_0.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_0.a_inv = "false";
defparam carry_13_ADD_0.PCK_LOCATION = "C18R21.lp0.add2.add0";
ADD1_A carry_9_ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[3]|qx_net  ),
	. ci ( \carry_9_ADD_2|co_net  ),
	. co ( \carry_9_ADD_3|co_net  ),
	. s ( \carry_9_ADD_3|s_net  )
);
defparam carry_9_ADD_3.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_3.a_inv = "true";
defparam carry_9_ADD_3.PCK_LOCATION = "C16R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[27]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .PCK_LOCATION = "C8R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[27] .always_en = 1;
REG glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg|qx_net  ),
	. di ( \ii3314|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_sec_vs_delay_flag_reg.always_en = 1;
LUT6 ii2421 (
	. xy ( \ii2421|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[5]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[4]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[3]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[2]|qx_net  )
);
defparam ii2421.PLACE_LOCATION = "C20R4.le_tile.le_guts.lp0.lut_0";
defparam ii2421.PCK_LOCATION = "C20R4.lp0.lut_0";
defparam ii2421.config_data = 64'b0000000000000010000000000000001000000000000000100000000000000010;
ADD1_A carry_13_ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1]|qx_net  ),
	. ci ( \carry_13_ADD_0|co_net  ),
	. co ( \carry_13_ADD_1|co_net  ),
	. s ( \carry_13_ADD_1|s_net  )
);
defparam carry_13_ADD_1.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_1.a_inv = "false";
defparam carry_13_ADD_1.PCK_LOCATION = "C18R21.lp0.add2.add0";
ADD1_A carry_9_ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[4]|qx_net  ),
	. ci ( \carry_9_ADD_3|co_net  ),
	. co ( \carry_9_ADD_4|co_net  ),
	. s ( \carry_9_ADD_4|s_net  )
);
defparam carry_9_ADD_4.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_4.a_inv = "true";
defparam carry_9_ADD_4.PCK_LOCATION = "C16R7.lp0.add2.add0";
LUT6 ii2422 (
	. xy ( \ii2422|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[1]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[11]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[10]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_sc1_rst_cnt_reg[0]|qx_net  ),
	. f1 ( \ii2421|xy_net  ),
	. f0 ( \ii2420|xy_net  )
);
defparam ii2422.PLACE_LOCATION = "C20R5.le_tile.le_guts.lp0.lut_0";
defparam ii2422.PCK_LOCATION = "C20R5.lp0.lut_0";
defparam ii2422.config_data = 64'b1111111111111111111111111111011111111111111111111111111111111111;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[28]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf.PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf.PCK_LOCATION = "C6R12.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .PLACE_LOCATION = "C10R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .PCK_LOCATION = "C10R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t11_reg_reg[2] .always_en = 1;
ADD1_A carry_13_ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2]|qx_net  ),
	. ci ( \carry_13_ADD_1|co_net  ),
	. co ( \carry_13_ADD_2|co_net  ),
	. s ( \carry_13_ADD_2|s_net  )
);
defparam carry_13_ADD_2.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_2.a_inv = "false";
defparam carry_13_ADD_2.PCK_LOCATION = "C18R21.lp0.add2.add0";
ADD1_A carry_9_ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[5]|qx_net  ),
	. ci ( \carry_9_ADD_4|co_net  ),
	. co ( \carry_9_ADD_5|co_net  ),
	. s ( \carry_9_ADD_5|s_net  )
);
defparam carry_9_ADD_5.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_5.a_inv = "true";
defparam carry_9_ADD_5.PCK_LOCATION = "C16R7.lp0.add2.add0";
LUT6 ii2423 (
	. xy ( \ii2423|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_fifo_sync_readen_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|dout[0]_net  )
);
defparam ii2423.PLACE_LOCATION = "C14R16.le_tile.le_guts.lp0.lut_0";
defparam ii2423.PCK_LOCATION = "C14R16.lp0.lut_0";
defparam ii2423.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62]|qx_net  ),
	. di ( \ii2214|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .PCK_LOCATION = "C16R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[62] .always_en = 0;
ADD1_A carry_13_ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3]|qx_net  ),
	. ci ( \carry_13_ADD_2|co_net  ),
	. co ( \carry_13_ADD_3|co_net  ),
	. s ( \carry_13_ADD_3|s_net  )
);
defparam carry_13_ADD_3.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_3.a_inv = "false";
defparam carry_13_ADD_3.PCK_LOCATION = "C18R21.lp0.add2.add0";
ADD1_A carry_9_ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[6]|qx_net  ),
	. ci ( \carry_9_ADD_5|co_net  ),
	. co ( \carry_9_ADD_6|co_net  ),
	. s ( \carry_9_ADD_6|s_net  )
);
defparam carry_9_ADD_6.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_6.a_inv = "true";
defparam carry_9_ADD_6.PCK_LOCATION = "C16R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_11__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[1] .always_en = 1;
LUT6 ii2424 (
	. xy ( \ii2424|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_fifo_sync_readen_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_fifo_sync_inst_u_inst|dout[1]_net  )
);
defparam ii2424.PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.lut_0";
defparam ii2424.PCK_LOCATION = "C16R15.lp0.lut_0";
defparam ii2424.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
ADD1_A carry_13_ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4]|qx_net  ),
	. ci ( \carry_13_ADD_3|co_net  ),
	. co ( \carry_13_ADD_4|co_net  ),
	. s ( \carry_13_ADD_4|s_net  )
);
defparam carry_13_ADD_4.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_4.a_inv = "false";
defparam carry_13_ADD_4.PCK_LOCATION = "C18R21.lp0.add2.add0";
ADD1_A carry_9_ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t2_out1_reg[7]|qx_net  ),
	. ci ( \carry_9_ADD_6|co_net  ),
	. co ( \carry_9_ADD_7|co_net  ),
	. s ( \carry_9_ADD_7|s_net  )
);
defparam carry_9_ADD_7.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_7.a_inv = "true";
defparam carry_9_ADD_7.PCK_LOCATION = "C16R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .PLACE_LOCATION = "C8R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .PCK_LOCATION = "C8R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[0] .always_en = 1;
LUT6 ii2425 (
	. xy ( \ii2425|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_rx_cmd_valid_dual_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[0]|qx_net  )
);
defparam ii2425.PLACE_LOCATION = "C4R8.le_tile.le_guts.lp0.lut_0";
defparam ii2425.PCK_LOCATION = "C4R8.lp0.lut_0";
defparam ii2425.config_data = 64'b0100000000000000000000000000000000000000000000000000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_data_process_frame_start_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0] .always_en = 1;
ADD1_A carry_13_ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5]|qx_net  ),
	. ci ( \carry_13_ADD_4|co_net  ),
	. co ( \carry_13_ADD_5|co_net  ),
	. s ( \carry_13_ADD_5|s_net  )
);
defparam carry_13_ADD_5.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_5.a_inv = "false";
defparam carry_13_ADD_5.PCK_LOCATION = "C18R21.lp0.add2.add0";
ADD1_A carry_9_ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_ADD_7|co_net  ),
	. co ( \carry_9_ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_ADD_8.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_ADD_8.a_inv = "false";
defparam carry_9_ADD_8.PCK_LOCATION = "C16R8.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_reg_reg_2_[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .PCK_LOCATION = "C18R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_In1p_reg[5] .always_en = 1;
LUT6 ii2426 (
	. xy ( \ii2426|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_cmd_dual_reg[5]|qx_net  ),
	. f0 ( \ii2425|xy_net  )
);
defparam ii2426.PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.lut_0";
defparam ii2426.PCK_LOCATION = "C6R6.lp0.lut_0";
defparam ii2426.config_data = 64'b1000111110001000100011111000100010001111100010001000111110001000;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[6]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[6]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7]|qx_net  ),
	. di ( \ii2502|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_6_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11]|qx_net  ),
	. di ( \ii2329|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .PCK_LOCATION = "C10R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11] .always_en = 0;
ADD1_A carry_13_ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6]|qx_net  ),
	. ci ( \carry_13_ADD_5|co_net  ),
	. co ( \carry_13_ADD_6|co_net  ),
	. s ( \carry_13_ADD_6|s_net  )
);
defparam carry_13_ADD_6.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_6.a_inv = "false";
defparam carry_13_ADD_6.PCK_LOCATION = "C18R21.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_12__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[4] .always_en = 1;
LUT6 ii2427 (
	. xy ( \ii2427|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_payload_valid_d_reg|qx_net  )
);
defparam ii2427.PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.lut_0";
defparam ii2427.PCK_LOCATION = "C10R7.lp0.lut_0";
defparam ii2427.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[4] .always_en = 1;
ADD1_A carry_13_ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7]|qx_net  ),
	. ci ( \carry_13_ADD_6|co_net  ),
	. co ( \carry_13_ADD_7|co_net  ),
	. s ( \carry_13_ADD_7|s_net  )
);
defparam carry_13_ADD_7.PLACE_LOCATION = "C18R21.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_7.a_inv = "false";
defparam carry_13_ADD_7.PCK_LOCATION = "C18R21.lp0.add2.add0";
LUT6 ii2428 (
	. xy ( \ii2428|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_data_process_first_3e_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_d_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  )
);
defparam ii2428.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.lut_0";
defparam ii2428.PCK_LOCATION = "C8R5.lp0.lut_0";
defparam ii2428.config_data = 64'b0101010100010000010101010001000001010101000100000101010100010000;
ADD1_A carry_13_ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8]|qx_net  ),
	. ci ( \carry_13_ADD_7|co_net  ),
	. co ( \carry_13_ADD_8|co_net  ),
	. s ( \carry_13_ADD_8|s_net  )
);
defparam carry_13_ADD_8.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_8.a_inv = "false";
defparam carry_13_ADD_8.PCK_LOCATION = "C18R22.lp0.add2.add0";
LUT6 ii2429 (
	. xy ( \ii2429|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_data_process_frame_start_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_data_process_first_3e_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_rx_hsync_reg|qx_net  )
);
defparam ii2429.PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.lut_0";
defparam ii2429.PCK_LOCATION = "C14R10.lp0.lut_0";
defparam ii2429.config_data = 64'b0011001100100000001100110010000000110011001000000011001100100000;
LUT6 ii2430 (
	. xy ( \ii2430|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t99_out1_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t105_out1_reg|qx_net  )
);
defparam ii2430.PLACE_LOCATION = "C20R26.le_tile.le_guts.lp0.lut_0";
defparam ii2430.PCK_LOCATION = "C20R26.lp0.lut_0";
defparam ii2430.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5]|qx_net  ),
	. di ( \ii2563|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5] .always_en = 1;
ADD1_A carry_13_ADD_9 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9]|qx_net  ),
	. ci ( \carry_13_ADD_8|co_net  ),
	. co ( \carry_13_ADD_9|co_net  ),
	. s ( \carry_13_ADD_9|s_net  )
);
defparam carry_13_ADD_9.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_13_ADD_9.a_inv = "false";
defparam carry_13_ADD_9.PCK_LOCATION = "C18R22.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[28]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[28] .always_en = 1;
LUT6 ii2431 (
	. xy ( \ii2431|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2431.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii2431.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii2431.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2432 (
	. xy ( \ii2432|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2432.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii2432.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii2432.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2433 (
	. xy ( \ii2433|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2433.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii2433.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii2433.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63]|qx_net  ),
	. di ( \ii2215|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2153|xy_net  ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .PLACE_LOCATION = "C16R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .PCK_LOCATION = "C16R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_cmd_byte_count_reg[63] .always_en = 0;
ADD1_A carry_8_ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_8_ADD_0|co_net  ),
	. s ( )
);
defparam carry_8_ADD_0.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_0.a_inv = "false";
defparam carry_8_ADD_0.PCK_LOCATION = "C14R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_11__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .PCK_LOCATION = "C18R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[2] .always_en = 1;
LUT6 ii2434 (
	. xy ( \ii2434|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2434.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii2434.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii2434.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_8_ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[1]|qx_net  ),
	. ci ( \carry_8_ADD_0|co_net  ),
	. co ( \carry_8_ADD_1|co_net  ),
	. s ( \carry_8_ADD_1|s_net  )
);
defparam carry_8_ADD_1.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_1.a_inv = "false";
defparam carry_8_ADD_1.PCK_LOCATION = "C14R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .PLACE_LOCATION = "C10R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .PCK_LOCATION = "C10R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[1] .always_en = 1;
LUT6 ii2435 (
	. xy ( \ii2435|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2435.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii2435.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii2435.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1] .always_en = 1;
ADD1_A carry_8_ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[2]|qx_net  ),
	. ci ( \carry_8_ADD_1|co_net  ),
	. co ( \carry_8_ADD_2|co_net  ),
	. s ( \carry_8_ADD_2|s_net  )
);
defparam carry_8_ADD_2.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_2.a_inv = "false";
defparam carry_8_ADD_2.PCK_LOCATION = "C14R17.lp0.add2.add0";
LUT6 ii2436 (
	. xy ( \ii2436|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2436.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2436.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2436.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[7]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[7]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[7] .always_en = 1;
ADD1_A carry_12_ADD_0 (
	. a ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_12_ADD_0|co_net  ),
	. s ( )
);
defparam carry_12_ADD_0.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_0.a_inv = "false";
defparam carry_12_ADD_0.PCK_LOCATION = "C14R22.lp0.add2.add0";
ADD1_A carry_8_ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[3]|qx_net  ),
	. ci ( \carry_8_ADD_2|co_net  ),
	. co ( \carry_8_ADD_3|co_net  ),
	. s ( \carry_8_ADD_3|s_net  )
);
defparam carry_8_ADD_3.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_3.a_inv = "false";
defparam carry_8_ADD_3.PCK_LOCATION = "C14R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_12__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[5] .always_en = 1;
LUT6 ii2437 (
	. xy ( \ii2437|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2437.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2437.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2437.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[5] .always_en = 1;
ADD1_A carry_12_ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[1]|qx_net  ),
	. ci ( \carry_12_ADD_0|co_net  ),
	. co ( \carry_12_ADD_1|co_net  ),
	. s ( \carry_12_ADD_1|s_net  )
);
defparam carry_12_ADD_1.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_1.a_inv = "false";
defparam carry_12_ADD_1.PCK_LOCATION = "C14R22.lp0.add2.add0";
ADD1_A carry_8_ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[4]|qx_net  ),
	. ci ( \carry_8_ADD_3|co_net  ),
	. co ( \carry_8_ADD_4|co_net  ),
	. s ( \carry_8_ADD_4|s_net  )
);
defparam carry_8_ADD_4.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_4.a_inv = "false";
defparam carry_8_ADD_4.PCK_LOCATION = "C14R17.lp0.add2.add0";
LUT6 ii2438 (
	. xy ( \ii2438|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_8_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2438.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2438.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2438.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
ADD1_A carry_12_ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[2]|qx_net  ),
	. ci ( \carry_12_ADD_1|co_net  ),
	. co ( \carry_12_ADD_2|co_net  ),
	. s ( \carry_12_ADD_2|s_net  )
);
defparam carry_12_ADD_2.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_2.a_inv = "false";
defparam carry_12_ADD_2.PCK_LOCATION = "C14R22.lp0.add2.add0";
ADD1_A carry_8_ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[5]|qx_net  ),
	. ci ( \carry_8_ADD_4|co_net  ),
	. co ( \carry_8_ADD_5|co_net  ),
	. s ( \carry_8_ADD_5|s_net  )
);
defparam carry_8_ADD_5.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_5.a_inv = "false";
defparam carry_8_ADD_5.PCK_LOCATION = "C14R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[0] .always_en = 1;
LUT6 ii2439 (
	. xy ( \ii2439|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2439.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2439.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2439.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2440 (
	. xy ( \ii2440|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2440.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2440.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2440.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6]|qx_net  ),
	. di ( \ii2564|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6] .always_en = 1;
ADD1_A carry_12_ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[3]|qx_net  ),
	. ci ( \carry_12_ADD_2|co_net  ),
	. co ( \carry_12_ADD_3|co_net  ),
	. s ( \carry_12_ADD_3|s_net  )
);
defparam carry_12_ADD_3.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_3.a_inv = "false";
defparam carry_12_ADD_3.PCK_LOCATION = "C14R22.lp0.add2.add0";
ADD1_A carry_8_ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[6]|qx_net  ),
	. ci ( \carry_8_ADD_5|co_net  ),
	. co ( \carry_8_ADD_6|co_net  ),
	. s ( \carry_8_ADD_6|s_net  )
);
defparam carry_8_ADD_6.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_6.a_inv = "false";
defparam carry_8_ADD_6.PCK_LOCATION = "C14R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[29]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[29] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[30]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[30] .always_en = 1;
LUT6 ii2441 (
	. xy ( \ii2441|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2441.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2441.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2441.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_12_ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[4]|qx_net  ),
	. ci ( \carry_12_ADD_3|co_net  ),
	. co ( \carry_12_ADD_4|co_net  ),
	. s ( \carry_12_ADD_4|s_net  )
);
defparam carry_12_ADD_4.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_4.a_inv = "false";
defparam carry_12_ADD_4.PCK_LOCATION = "C14R22.lp0.add2.add0";
ADD1_A carry_8_ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_sync_delay_hcnt_reg[7]|qx_net  ),
	. ci ( \carry_8_ADD_6|co_net  ),
	. co ( ),
	. s ( \carry_8_ADD_7|s_net  )
);
defparam carry_8_ADD_7.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_8_ADD_7.a_inv = "false";
defparam carry_8_ADD_7.PCK_LOCATION = "C14R17.lp0.add2.add0";
LUT6 ii2442 (
	. xy ( \ii2442|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2442.PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.lut_0";
defparam ii2442.PCK_LOCATION = "C20R10.lp0.lut_0";
defparam ii2442.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_12_ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[5]|qx_net  ),
	. ci ( \carry_12_ADD_4|co_net  ),
	. co ( \carry_12_ADD_5|co_net  ),
	. s ( \carry_12_ADD_5|s_net  )
);
defparam carry_12_ADD_5.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_5.a_inv = "false";
defparam carry_12_ADD_5.PCK_LOCATION = "C14R22.lp0.add2.add0";
LUT6 ii2443 (
	. xy ( \ii2443|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2443.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2443.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2443.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_12_ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[6]|qx_net  ),
	. ci ( \carry_12_ADD_5|co_net  ),
	. co ( \carry_12_ADD_6|co_net  ),
	. s ( \carry_12_ADD_6|s_net  )
);
defparam carry_12_ADD_6.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_6.a_inv = "false";
defparam carry_12_ADD_6.PCK_LOCATION = "C14R22.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_11__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[3] .always_en = 1;
LUT6 ii2444 (
	. xy ( \ii2444|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2444.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2444.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2444.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_12_ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[7]|qx_net  ),
	. ci ( \carry_12_ADD_6|co_net  ),
	. co ( \carry_12_ADD_7|co_net  ),
	. s ( \carry_12_ADD_7|s_net  )
);
defparam carry_12_ADD_7.PLACE_LOCATION = "C14R22.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_7.a_inv = "false";
defparam carry_12_ADD_7.PCK_LOCATION = "C14R22.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .PCK_LOCATION = "C14R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[2] .always_en = 1;
LUT6 ii2445 (
	. xy ( \ii2445|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2445.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2445.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2445.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
ADD1_A carry_12_ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[8]|qx_net  ),
	. ci ( \carry_12_ADD_7|co_net  ),
	. co ( \carry_12_ADD_8|co_net  ),
	. s ( \carry_12_ADD_8|s_net  )
);
defparam carry_12_ADD_8.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_8.a_inv = "false";
defparam carry_12_ADD_8.PCK_LOCATION = "C14R23.lp0.add2.add0";
LUT6 ii2446 (
	. xy ( \ii2446|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2446.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2446.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2446.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[8]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[8]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[8] .always_en = 1;
ADD1_A carry_12_ADD_9 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_tx_line_cnt_reg[9]|qx_net  ),
	. ci ( \carry_12_ADD_8|co_net  ),
	. co ( \carry_12_ADD_9|co_net  ),
	. s ( \carry_12_ADD_9|s_net  )
);
defparam carry_12_ADD_9.PLACE_LOCATION = "C14R23.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_ADD_9.a_inv = "false";
defparam carry_12_ADD_9.PCK_LOCATION = "C14R23.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_12__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[6] .always_en = 1;
LUT6 ii2447 (
	. xy ( \ii2447|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2447.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.lut_0";
defparam ii2447.PCK_LOCATION = "C16R17.lp0.lut_0";
defparam ii2447.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[18]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf.PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf.PCK_LOCATION = "C16R15.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[6] .always_en = 1;
LUT6 ii2448 (
	. xy ( \ii2448|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2448.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.lut_0";
defparam ii2448.PCK_LOCATION = "C16R17.lp0.lut_0";
defparam ii2448.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[1] .always_en = 1;
LUT6 ii2449 (
	. xy ( \ii2449|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2449.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.lut_0";
defparam ii2449.PCK_LOCATION = "C16R17.lp0.lut_0";
defparam ii2449.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2450 (
	. xy ( \ii2450|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2450.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.lut_0";
defparam ii2450.PCK_LOCATION = "C16R17.lp0.lut_0";
defparam ii2450.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
FIFO9K mcu_arbiter_u_pfifo_u_inst (
	. dout ( {
		/* dout [31] */ \mcu_arbiter_u_pfifo_u_inst|dout[31]_net ,
		/* dout [30] */ \mcu_arbiter_u_pfifo_u_inst|dout[30]_net ,
		/* dout [29] */ \mcu_arbiter_u_pfifo_u_inst|dout[29]_net ,
		/* dout [28] */ \mcu_arbiter_u_pfifo_u_inst|dout[28]_net ,
		/* dout [27] */ \mcu_arbiter_u_pfifo_u_inst|dout[27]_net ,
		/* dout [26] */ \mcu_arbiter_u_pfifo_u_inst|dout[26]_net ,
		/* dout [25] */ \mcu_arbiter_u_pfifo_u_inst|dout[25]_net ,
		/* dout [24] */ \mcu_arbiter_u_pfifo_u_inst|dout[24]_net ,
		/* dout [23] */ \mcu_arbiter_u_pfifo_u_inst|dout[23]_net ,
		/* dout [22] */ \mcu_arbiter_u_pfifo_u_inst|dout[22]_net ,
		/* dout [21] */ \mcu_arbiter_u_pfifo_u_inst|dout[21]_net ,
		/* dout [20] */ \mcu_arbiter_u_pfifo_u_inst|dout[20]_net ,
		/* dout [19] */ \mcu_arbiter_u_pfifo_u_inst|dout[19]_net ,
		/* dout [18] */ \mcu_arbiter_u_pfifo_u_inst|dout[18]_net ,
		/* dout [17] */ \mcu_arbiter_u_pfifo_u_inst|dout[17]_net ,
		/* dout [16] */ \mcu_arbiter_u_pfifo_u_inst|dout[16]_net ,
		/* dout [15] */ \mcu_arbiter_u_pfifo_u_inst|dout[15]_net ,
		/* dout [14] */ \mcu_arbiter_u_pfifo_u_inst|dout[14]_net ,
		/* dout [13] */ \mcu_arbiter_u_pfifo_u_inst|dout[13]_net ,
		/* dout [12] */ \mcu_arbiter_u_pfifo_u_inst|dout[12]_net ,
		/* dout [11] */ \mcu_arbiter_u_pfifo_u_inst|dout[11]_net ,
		/* dout [10] */ \mcu_arbiter_u_pfifo_u_inst|dout[10]_net ,
		/* dout [9] */ \mcu_arbiter_u_pfifo_u_inst|dout[9]_net ,
		/* dout [8] */ \mcu_arbiter_u_pfifo_u_inst|dout[8]_net ,
		/* dout [7] */ \mcu_arbiter_u_pfifo_u_inst|dout[7]_net ,
		/* dout [6] */ \mcu_arbiter_u_pfifo_u_inst|dout[6]_net ,
		/* dout [5] */ \mcu_arbiter_u_pfifo_u_inst|dout[5]_net ,
		/* dout [4] */ \mcu_arbiter_u_pfifo_u_inst|dout[4]_net ,
		/* dout [3] */ \mcu_arbiter_u_pfifo_u_inst|dout[3]_net ,
		/* dout [2] */ \mcu_arbiter_u_pfifo_u_inst|dout[2]_net ,
		/* dout [1] */ \mcu_arbiter_u_pfifo_u_inst|dout[1]_net ,
		/* dout [0] */ \mcu_arbiter_u_pfifo_u_inst|dout[0]_net 
	} ),
	. doutp ( )
,
	. din ( {
		/* din [31] */ \GND_0_inst|Y_net ,
		/* din [30] */ \GND_0_inst|Y_net ,
		/* din [29] */ \GND_0_inst|Y_net ,
		/* din [28] */ \GND_0_inst|Y_net ,
		/* din [27] */ \GND_0_inst|Y_net ,
		/* din [26] */ \GND_0_inst|Y_net ,
		/* din [25] */ \GND_0_inst|Y_net ,
		/* din [24] */ \GND_0_inst|Y_net ,
		/* din [23] */ \GND_0_inst|Y_net ,
		/* din [22] */ \GND_0_inst|Y_net ,
		/* din [21] */ \GND_0_inst|Y_net ,
		/* din [20] */ \GND_0_inst|Y_net ,
		/* din [19] */ \GND_0_inst|Y_net ,
		/* din [18] */ \GND_0_inst|Y_net ,
		/* din [17] */ \GND_0_inst|Y_net ,
		/* din [16] */ \GND_0_inst|Y_net ,
		/* din [15] */ \GND_0_inst|Y_net ,
		/* din [14] */ \GND_0_inst|Y_net ,
		/* din [13] */ \GND_0_inst|Y_net ,
		/* din [12] */ \GND_0_inst|Y_net ,
		/* din [11] */ \GND_0_inst|Y_net ,
		/* din [10] */ \GND_0_inst|Y_net ,
		/* din [9] */ \GND_0_inst|Y_net ,
		/* din [8] */ \GND_0_inst|Y_net ,
		/* din [7] */ \u_8051_u_h6_8051|memdatao_comb[7]_net ,
		/* din [6] */ \u_8051_u_h6_8051|memdatao_comb[6]_net ,
		/* din [5] */ \u_8051_u_h6_8051|memdatao_comb[5]_net ,
		/* din [4] */ \u_8051_u_h6_8051|memdatao_comb[4]_net ,
		/* din [3] */ \u_8051_u_h6_8051|memdatao_comb[3]_net ,
		/* din [2] */ \u_8051_u_h6_8051|memdatao_comb[2]_net ,
		/* din [1] */ \u_8051_u_h6_8051|memdatao_comb[1]_net ,
		/* din [0] */ \u_8051_u_h6_8051|memdatao_comb[0]_net 
	} ),
	. dinp ( {
		/* dinp [3] */ \GND_0_inst|Y_net ,
		/* dinp [2] */ \GND_0_inst|Y_net ,
		/* dinp [1] */ \GND_0_inst|Y_net ,
		/* dinp [0] (nc) */ nc568 
	} ),
	. writeclk ( \u_pll_pll_u0|CO3_net  ),
	. readclk ( \u_gbuf_u_gbuf|out_net  ),
	. writeen ( \ii2040|xy_net  ),
	. readen ( \ii2036|xy_net  ),
	. reset ( \ii2037|xy_net  ),
	. regce ( ),
	. writesave ( \GND_0_inst|Y_net  ),
	. writedrop ( \GND_0_inst|Y_net  ),
	. full ( ),
	. empty ( ),
	. almostfull ( ),
	. almostempty ( ),
	. overflow ( ),
	. underflow ( ),
	. writedropflag ( )
);
defparam mcu_arbiter_u_pfifo_u_inst.readwidth = 36;
defparam mcu_arbiter_u_pfifo_u_inst.PLACE_LOCATION = "C12R29.emb_guts.u0_emb_top.emb18k_wrapper.u0_emb18k_core.bram9k_0";
defparam mcu_arbiter_u_pfifo_u_inst.use_parity = 0;
defparam mcu_arbiter_u_pfifo_u_inst.writeclk_inv = 0;
defparam mcu_arbiter_u_pfifo_u_inst.peek = 0;
defparam mcu_arbiter_u_pfifo_u_inst.PCK_LOCATION = "C12R29.u0_emb_top.emb18k_wrapper.u0_emb18k_core.bram9k_0";
defparam mcu_arbiter_u_pfifo_u_inst.readclk_inv = 0;
defparam mcu_arbiter_u_pfifo_u_inst.outreg = 0;
defparam mcu_arbiter_u_pfifo_u_inst.writewidth = 9;
defparam mcu_arbiter_u_pfifo_u_inst.almostfullth = 8;
defparam mcu_arbiter_u_pfifo_u_inst.almostemptyth = 6;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7]|qx_net  ),
	. di ( \ii2565|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[31]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .PCK_LOCATION = "C16R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[31] .always_en = 1;
LUT6 ii2451 (
	. xy ( \ii2451|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2451.PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.lut_0";
defparam ii2451.PCK_LOCATION = "C16R17.lp0.lut_0";
defparam ii2451.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2452 (
	. xy ( \ii2452|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2452.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2452.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2452.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2453 (
	. xy ( \ii2453|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2453.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2453.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2453.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
ADD1_A carry_11_ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \GND_0_inst|Y_net  ),
	. co ( \carry_11_ADD_0|co_net  ),
	. s ( )
);
defparam carry_11_ADD_0.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_0.a_inv = "false";
defparam carry_11_ADD_0.PCK_LOCATION = "C18R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_11__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[4] .always_en = 1;
LUT6 ii2454 (
	. xy ( \ii2454|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2454.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2454.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2454.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
ADD1_A carry_11_ADD_1 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[1]|qx_net  ),
	. ci ( \carry_11_ADD_0|co_net  ),
	. co ( \carry_11_ADD_1|co_net  ),
	. s ( \carry_11_ADD_1|s_net  )
);
defparam carry_11_ADD_1.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_1.a_inv = "false";
defparam carry_11_ADD_1.PCK_LOCATION = "C18R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .PCK_LOCATION = "C16R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[3] .always_en = 1;
LUT6 ii2455 (
	. xy ( \ii2455|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2455.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2455.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2455.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_11_ADD_2 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2]|qx_net  ),
	. ci ( \carry_11_ADD_1|co_net  ),
	. co ( \carry_11_ADD_2|co_net  ),
	. s ( \carry_11_ADD_2|s_net  )
);
defparam carry_11_ADD_2.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_2.a_inv = "false";
defparam carry_11_ADD_2.PCK_LOCATION = "C18R17.lp0.add2.add0";
LUT6 ii2456 (
	. xy ( \ii2456|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2456.PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.lut_0";
defparam ii2456.PCK_LOCATION = "C18R16.lp0.lut_0";
defparam ii2456.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \uut_dataReadBack_mipi_periph_tx_payload_reg[9]  (
	. qx ( \uut_dataReadBack_mipi_periph_tx_payload_reg[9]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .latch_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .init = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .PLACE_LOCATION = "C6R3.le_tile.le_guts.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .sr_inv = 1;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .sync_mode = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .no_sr = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .sr_value = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .PCK_LOCATION = "C6R3.lp0.reg0";
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .clk_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .en_inv = 0;
defparam \uut_dataReadBack_mipi_periph_tx_payload_reg[9] .always_en = 1;
ADD1_A carry_11_ADD_3 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3]|qx_net  ),
	. ci ( \carry_11_ADD_2|co_net  ),
	. co ( \carry_11_ADD_3|co_net  ),
	. s ( \carry_11_ADD_3|s_net  )
);
defparam carry_11_ADD_3.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_3.a_inv = "false";
defparam carry_11_ADD_3.PCK_LOCATION = "C18R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_12__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[7] .always_en = 1;
LUT6 ii2457 (
	. xy ( \ii2457|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2457.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2457.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2457.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .PCK_LOCATION = "C14R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t101_out1_reg[7] .always_en = 1;
REG glue_rx_packet_tx_packet_fifo_empty_reg (
	. qx ( \glue_rx_packet_tx_packet_fifo_empty_reg|qx_net  ),
	. di ( \ii2139|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_fifo_empty_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.init = 0;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.PLACE_LOCATION = "C14R25.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_fifo_empty_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.sr_value = 1;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.PCK_LOCATION = "C14R25.lp0.reg0";
defparam glue_rx_packet_tx_packet_fifo_empty_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_fifo_empty_reg.always_en = 1;
ADD1_A carry_11_ADD_4 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4]|qx_net  ),
	. ci ( \carry_11_ADD_3|co_net  ),
	. co ( \carry_11_ADD_4|co_net  ),
	. s ( \carry_11_ADD_4|s_net  )
);
defparam carry_11_ADD_4.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_4.a_inv = "false";
defparam carry_11_ADD_4.PCK_LOCATION = "C18R17.lp0.add2.add0";
LUT6 ii2458 (
	. xy ( \ii2458|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2458.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2458.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2458.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_11_ADD_5 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5]|qx_net  ),
	. ci ( \carry_11_ADD_4|co_net  ),
	. co ( \carry_11_ADD_5|co_net  ),
	. s ( \carry_11_ADD_5|s_net  )
);
defparam carry_11_ADD_5.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_5.a_inv = "false";
defparam carry_11_ADD_5.PCK_LOCATION = "C18R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[2] .always_en = 1;
LUT6 ii2459 (
	. xy ( \ii2459|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2459.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2459.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2459.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2460 (
	. xy ( \ii2460|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2460.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2460.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2460.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8]|qx_net  ),
	. di ( \ii2566|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8] .always_en = 1;
ADD1_A carry_11_ADD_6 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6]|qx_net  ),
	. ci ( \carry_11_ADD_5|co_net  ),
	. co ( \carry_11_ADD_6|co_net  ),
	. s ( \carry_11_ADD_6|s_net  )
);
defparam carry_11_ADD_6.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_6.a_inv = "false";
defparam carry_11_ADD_6.PCK_LOCATION = "C18R17.lp0.add2.add0";
LUT6 ii2461 (
	. xy ( \ii2461|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2461.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2461.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2461.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
ADD1_A carry_11_ADD_7 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7]|qx_net  ),
	. ci ( \carry_11_ADD_6|co_net  ),
	. co ( \carry_11_ADD_7|co_net  ),
	. s ( \carry_11_ADD_7|s_net  )
);
defparam carry_11_ADD_7.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_7.a_inv = "false";
defparam carry_11_ADD_7.PCK_LOCATION = "C18R17.lp0.add2.add0";
LUT6 ii2462 (
	. xy ( \ii2462|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2462.PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.lut_0";
defparam ii2462.PCK_LOCATION = "C16R16.lp0.lut_0";
defparam ii2462.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .PLACE_LOCATION = "C6R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .PCK_LOCATION = "C6R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[0] .always_en = 1;
ADD1_A carry_11_ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8]|qx_net  ),
	. ci ( \carry_11_ADD_7|co_net  ),
	. co ( \carry_11_ADD_8|co_net  ),
	. s ( \carry_11_ADD_8|s_net  )
);
defparam carry_11_ADD_8.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_8.a_inv = "false";
defparam carry_11_ADD_8.PCK_LOCATION = "C18R18.lp0.add2.add0";
LUT6 ii2463 (
	. xy ( \ii2463|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2463.PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.lut_0";
defparam ii2463.PCK_LOCATION = "C8R6.lp0.lut_0";
defparam ii2463.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_11_ADD_9 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9]|qx_net  ),
	. ci ( \carry_11_ADD_8|co_net  ),
	. co ( \carry_11_ADD_9|co_net  ),
	. s ( \carry_11_ADD_9|s_net  )
);
defparam carry_11_ADD_9.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.add2.add0";
defparam carry_11_ADD_9.a_inv = "false";
defparam carry_11_ADD_9.PCK_LOCATION = "C18R18.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .PCK_LOCATION = "C14R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t7_out1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_11__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[5] .always_en = 1;
LUT6 ii2464 (
	. xy ( \ii2464|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2464.PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.lut_0";
defparam ii2464.PCK_LOCATION = "C8R6.lp0.lut_0";
defparam ii2464.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[4] .always_en = 1;
LUT6 ii2465 (
	. xy ( \ii2465|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2465.PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.lut_0";
defparam ii2465.PCK_LOCATION = "C8R6.lp0.lut_0";
defparam ii2465.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_9_6__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_6__ADD_0|co_net  ),
	. s ( \carry_9_6__ADD_0|s_net  )
);
defparam carry_9_6__ADD_0.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_0.a_inv = "true";
defparam carry_9_6__ADD_0.PCK_LOCATION = "C20R16.lp0.add2.add0";
LUT6 ii2466 (
	. xy ( \ii2466|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2466.PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.lut_0";
defparam ii2466.PCK_LOCATION = "C8R6.lp0.lut_0";
defparam ii2466.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_9_6__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1]|qx_net  ),
	. ci ( \carry_9_6__ADD_0|co_net  ),
	. co ( \carry_9_6__ADD_1|co_net  ),
	. s ( \carry_9_6__ADD_1|s_net  )
);
defparam carry_9_6__ADD_1.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_1.a_inv = "true";
defparam carry_9_6__ADD_1.PCK_LOCATION = "C20R16.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8]|qx_net  ),
	. di ( \ii2992|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In2p_reg[8] .always_en = 1;
LUT6 ii2467 (
	. xy ( \ii2467|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2467.PLACE_LOCATION = "C8R6.le_tile.le_guts.lp0.lut_0";
defparam ii2467.PCK_LOCATION = "C8R6.lp0.lut_0";
defparam ii2467.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[3] .always_en = 1;
ADD1_A carry_9_6__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2]|qx_net  ),
	. ci ( \carry_9_6__ADD_1|co_net  ),
	. co ( \carry_9_6__ADD_2|co_net  ),
	. s ( \carry_9_6__ADD_2|s_net  )
);
defparam carry_9_6__ADD_2.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_2.a_inv = "true";
defparam carry_9_6__ADD_2.PCK_LOCATION = "C20R16.lp0.add2.add0";
LUT6 ii2468 (
	. xy ( \ii2468|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2468.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2468.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2468.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_9_6__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[3]|qx_net  ),
	. ci ( \carry_9_6__ADD_2|co_net  ),
	. co ( \carry_9_6__ADD_3|co_net  ),
	. s ( \carry_9_6__ADD_3|s_net  )
);
defparam carry_9_6__ADD_3.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_3.a_inv = "true";
defparam carry_9_6__ADD_3.PCK_LOCATION = "C20R16.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[3] .always_en = 1;
LUT6 ii2469 (
	. xy ( \ii2469|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2469.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2469.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2469.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2470 (
	. xy ( \ii2470|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2470.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2470.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2470.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_1_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9]|qx_net  ),
	. di ( \ii2567|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .PCK_LOCATION = "C18R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9] .always_en = 1;
ADD1_A carry_9_6__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[4]|qx_net  ),
	. ci ( \carry_9_6__ADD_3|co_net  ),
	. co ( \carry_9_6__ADD_4|co_net  ),
	. s ( \carry_9_6__ADD_4|s_net  )
);
defparam carry_9_6__ADD_4.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_4.a_inv = "true";
defparam carry_9_6__ADD_4.PCK_LOCATION = "C20R16.lp0.add2.add0";
LUT6 ii2471 (
	. xy ( \ii2471|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2471.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2471.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2471.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_9_6__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[5]|qx_net  ),
	. ci ( \carry_9_6__ADD_4|co_net  ),
	. co ( \carry_9_6__ADD_5|co_net  ),
	. s ( \carry_9_6__ADD_5|s_net  )
);
defparam carry_9_6__ADD_5.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_5.a_inv = "true";
defparam carry_9_6__ADD_5.PCK_LOCATION = "C20R16.lp0.add2.add0";
LUT6 ii2472 (
	. xy ( \ii2472|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2472.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2472.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2472.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .PLACE_LOCATION = "C8R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .PCK_LOCATION = "C8R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[1] .always_en = 1;
ADD1_A carry_9_6__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[6]|qx_net  ),
	. ci ( \carry_9_6__ADD_5|co_net  ),
	. co ( \carry_9_6__ADD_6|co_net  ),
	. s ( \carry_9_6__ADD_6|s_net  )
);
defparam carry_9_6__ADD_6.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_6.a_inv = "true";
defparam carry_9_6__ADD_6.PCK_LOCATION = "C20R16.lp0.add2.add0";
LUT6 ii2473 (
	. xy ( \ii2473|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2473.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2473.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2473.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_9_6__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[7]|qx_net  ),
	. ci ( \carry_9_6__ADD_6|co_net  ),
	. co ( \carry_9_6__ADD_7|co_net  ),
	. s ( \carry_9_6__ADD_7|s_net  )
);
defparam carry_9_6__ADD_7.PLACE_LOCATION = "C20R16.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_7.a_inv = "true";
defparam carry_9_6__ADD_7.PCK_LOCATION = "C20R16.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_11__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[6] .always_en = 1;
LUT6 ii2474 (
	. xy ( \ii2474|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2474.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2474.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2474.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
ADD1_A carry_9_6__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_6__ADD_7|co_net  ),
	. co ( \carry_9_6__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_6__ADD_8.PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_6__ADD_8.a_inv = "false";
defparam carry_9_6__ADD_8.PCK_LOCATION = "C20R17.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[5] .always_en = 1;
LUT6 ii2475 (
	. xy ( \ii2475|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2475.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2475.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2475.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly (
	. xy ( \u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \u0_mipi1_clkdly_genblk1_2__u_mipi_clkdly|xy_net  )
);
defparam u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly.PLACE_LOCATION = "C20R23.le_tile.le_guts.lp0.lut_1";
defparam u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly.PCK_LOCATION = "NONE";
defparam u0_mipi1_clkdly_genblk1_1__u_mipi_clkdly.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2476 (
	. xy ( \ii2476|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2476.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2476.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2476.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[0] .always_en = 1;
LUT6 ii2477 (
	. xy ( \ii2477|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2477.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2477.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2477.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[4] .always_en = 1;
LUT6 ii2478 (
	. xy ( \ii2478|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2478.PLACE_LOCATION = "C8R7.le_tile.le_guts.lp0.lut_0";
defparam ii2478.PCK_LOCATION = "C8R7.lp0.lut_0";
defparam ii2478.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[4] .always_en = 1;
LUT6 ii2479 (
	. xy ( \ii2479|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2479.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2479.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2479.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2480 (
	. xy ( \ii2480|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2480.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2480.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2480.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2481 (
	. xy ( \ii2481|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2481.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.lut_0";
defparam ii2481.PCK_LOCATION = "C8R8.lp0.lut_0";
defparam ii2481.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2482 (
	. xy ( \ii2482|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2482.PLACE_LOCATION = "C8R8.le_tile.le_guts.lp0.lut_0";
defparam ii2482.PCK_LOCATION = "C8R8.lp0.lut_0";
defparam ii2482.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .PLACE_LOCATION = "C10R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .PCK_LOCATION = "C10R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[2] .always_en = 1;
LUT6 ii2483 (
	. xy ( \ii2483|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2483.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2483.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2483.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_11__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .PCK_LOCATION = "C20R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[7] .always_en = 1;
LUT6 ii2484 (
	. xy ( \ii2484|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2484.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2484.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2484.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[6] .always_en = 1;
LUT6 ii2485 (
	. xy ( \ii2485|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2485.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2485.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2485.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg|qx_net  ),
	. di ( \ii2426|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.PLACE_LOCATION = "C6R6.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.PCK_LOCATION = "C6R6.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_data_3Eh_valid_reg.always_en = 1;
LUT6 ii2486 (
	. xy ( \ii2486|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_2_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2486.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2486.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2486.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG glue_rx_packet_tx_packet_rx_vsync_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_vsync_reg|qx_net  ),
	. di ( \ii2295|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_vsync_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.PLACE_LOCATION = "C16R5.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_vsync_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.PCK_LOCATION = "C16R5.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_vsync_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_vsync_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t103_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .PLACE_LOCATION = "C20R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .PCK_LOCATION = "C20R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t4_out1_1_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[1] .always_en = 1;
LUT6 ii2487 (
	. xy ( \ii2487|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2487.PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.lut_0";
defparam ii2487.PCK_LOCATION = "C14R8.lp0.lut_0";
defparam ii2487.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[5] .always_en = 1;
LUT6 ii2488 (
	. xy ( \ii2488|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2488.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2488.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2488.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[5] .always_en = 1;
LUT6 ii2489 (
	. xy ( \ii2489|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2489.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2489.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2489.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2490 (
	. xy ( \ii2490|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2490.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2490.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2490.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2500 (
	. xy ( \ii2500|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2500.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2500.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2500.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2491 (
	. xy ( \ii2491|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2491.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2491.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2491.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2501 (
	. xy ( \ii2501|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2501.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2501.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2501.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2492 (
	. xy ( \ii2492|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2492.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2492.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2492.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2502 (
	. xy ( \ii2502|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2502.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2502.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2502.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_0_[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .PLACE_LOCATION = "C18R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .PCK_LOCATION = "C18R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_reg_reg_1_[3] .always_en = 1;
LUT6 ii2493 (
	. xy ( \ii2493|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2493.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2493.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2493.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2503 (
	. xy ( \ii2503|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2503.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2503.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2503.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8]|qx_net  ),
	. di ( \ii3282|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .PLACE_LOCATION = "C20R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .PCK_LOCATION = "C20R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In2p_reg[8] .always_en = 1;
LUT6 ii2494 (
	. xy ( \ii2494|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_3_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2494.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2494.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2494.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2504 (
	. xy ( \ii2504|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2504.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2504.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2504.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_12_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .PLACE_LOCATION = "C18R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .PCK_LOCATION = "C18R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In3p_reg[7] .always_en = 1;
LUT6 ii2495 (
	. xy ( \ii2495|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2495.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2495.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2495.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2505 (
	. xy ( \ii2505|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2505.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2505.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2505.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2496 (
	. xy ( \ii2496|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2496.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2496.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2496.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2506 (
	. xy ( \ii2506|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2506.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2506.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2506.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .PCK_LOCATION = "C16R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[2] .always_en = 1;
LUT6 ii2497 (
	. xy ( \ii2497|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2497.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2497.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2497.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2507 (
	. xy ( \ii2507|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2507.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2507.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2507.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[6] .always_en = 1;
LUT6 ii2498 (
	. xy ( \ii2498|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2498.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2498.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2498.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2508 (
	. xy ( \ii2508|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2508.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2508.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2508.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[6] .always_en = 1;
LUT6 ii2499 (
	. xy ( \ii2499|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2499.PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.lut_0";
defparam ii2499.PCK_LOCATION = "C20R19.lp0.lut_0";
defparam ii2499.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2509 (
	. xy ( \ii2509|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2509.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2509.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2509.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2510 (
	. xy ( \ii2510|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2510.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2510.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2510.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2511 (
	. xy ( \ii2511|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2511.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.lut_0";
defparam ii2511.PCK_LOCATION = "C18R14.lp0.lut_0";
defparam ii2511.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2512 (
	. xy ( \ii2512|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2512.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.lut_0";
defparam ii2512.PCK_LOCATION = "C18R14.lp0.lut_0";
defparam ii2512.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0] .always_en = 1;
LUT6 ii2513 (
	. xy ( \ii2513|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2513.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.lut_0";
defparam ii2513.PCK_LOCATION = "C18R14.lp0.lut_0";
defparam ii2513.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2514 (
	. xy ( \ii2514|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2514.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii2514.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii2514.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2515 (
	. xy ( \ii2515|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2515.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii2515.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii2515.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2516 (
	. xy ( \ii2516|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2516.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii2516.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii2516.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0]|qx_net  ),
	. di ( \ii2487|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[3] .always_en = 1;
LUT6 ii2517 (
	. xy ( \ii2517|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2517.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii2517.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii2517.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .PLACE_LOCATION = "C16R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .PCK_LOCATION = "C16R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[7] .always_en = 1;
LUT6 ii2518 (
	. xy ( \ii2518|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2518.PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.lut_0";
defparam ii2518.PCK_LOCATION = "C20R14.lp0.lut_0";
defparam ii2518.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .PCK_LOCATION = "C16R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[7] .always_en = 1;
LUT6 ii2519 (
	. xy ( \ii2519|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[4]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2519.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.lut_0";
defparam ii2519.PCK_LOCATION = "C18R14.lp0.lut_0";
defparam ii2519.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2520 (
	. xy ( \ii2520|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[5]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2520.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.lut_0";
defparam ii2520.PCK_LOCATION = "C18R14.lp0.lut_0";
defparam ii2520.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. di ( \ii2617|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .PLACE_LOCATION = "C8R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .PCK_LOCATION = "C8R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10] .always_en = 1;
LUT6 ii2521 (
	. xy ( \ii2521|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[6]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2521.PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.lut_0";
defparam ii2521.PCK_LOCATION = "C18R14.lp0.lut_0";
defparam ii2521.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2522 (
	. xy ( \ii2522|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[7]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2522.PLACE_LOCATION = "C18R13.le_tile.le_guts.lp0.lut_0";
defparam ii2522.PCK_LOCATION = "C18R13.lp0.lut_0";
defparam ii2522.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1] .always_en = 1;
LUT6 ii2523 (
	. xy ( \ii2523|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[8]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2523.PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.lut_0";
defparam ii2523.PCK_LOCATION = "C20R13.lp0.lut_0";
defparam ii2523.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[14]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .PLACE_LOCATION = "C20R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .PCK_LOCATION = "C20R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[0] .always_en = 1;
LUT6 ii2524 (
	. xy ( \ii2524|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[9]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  )
);
defparam ii2524.PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.lut_0";
defparam ii2524.PCK_LOCATION = "C20R13.lp0.lut_0";
defparam ii2524.config_data = 64'b0000000011111111000000001111111000000000111111110000000011111110;
LUT6 ii2525 (
	. xy ( \ii2525|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[10]_net  )
);
defparam ii2525.PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.lut_0";
defparam ii2525.PCK_LOCATION = "C20R13.lp0.lut_0";
defparam ii2525.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
LUT6 ii2526 (
	. xy ( \ii2526|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[15]_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[14]_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[13]_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[12]_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_7_i73_mac_u0|a_mac_out[11]_net  )
);
defparam ii2526.PLACE_LOCATION = "C20R13.le_tile.le_guts.lp0.lut_0";
defparam ii2526.PCK_LOCATION = "C20R13.lp0.lut_0";
defparam ii2526.config_data = 64'b0000000000000000111111111111111000000000000000001111111111111110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1]|qx_net  ),
	. di ( \ii2488|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[4] .always_en = 1;
REG mcu_arbiter_fifo_clr_f_reg (
	. qx ( \mcu_arbiter_fifo_clr_f_reg|qx_net  ),
	. di ( \mcu_arbiter_func_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_fifo_clr_f_reg.latch_mode = 0;
defparam mcu_arbiter_fifo_clr_f_reg.init = 0;
defparam mcu_arbiter_fifo_clr_f_reg.PLACE_LOCATION = "C4R19.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_fifo_clr_f_reg.sr_inv = 1;
defparam mcu_arbiter_fifo_clr_f_reg.sync_mode = 0;
defparam mcu_arbiter_fifo_clr_f_reg.no_sr = 0;
defparam mcu_arbiter_fifo_clr_f_reg.sr_value = 0;
defparam mcu_arbiter_fifo_clr_f_reg.PCK_LOCATION = "C4R19.lp0.reg0";
defparam mcu_arbiter_fifo_clr_f_reg.clk_inv = 0;
defparam mcu_arbiter_fifo_clr_f_reg.en_inv = 0;
defparam mcu_arbiter_fifo_clr_f_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[10] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8]|qx_net  ),
	. di ( \ii2963|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .PLACE_LOCATION = "C10R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .PCK_LOCATION = "C10R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In2p_reg[8] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. di ( \ii2621|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[15]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .PLACE_LOCATION = "C20R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .PCK_LOCATION = "C20R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2]|qx_net  ),
	. di ( \ii2489|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t34_out1_1_reg[9] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[11]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[11] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. di ( \ii2625|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[16]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .PLACE_LOCATION = "C20R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .PCK_LOCATION = "C20R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3]|qx_net  ),
	. di ( \ii2490|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[6] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[12]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[12] .always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0]|qx_net  ),
	. di ( \ii2296|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[0] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. di ( \ii2629|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[17]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .PLACE_LOCATION = "C20R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .PCK_LOCATION = "C20R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[3] .always_en = 1;
LUT6 ii2555 (
	. xy ( \ii2555|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  )
);
defparam ii2555.PLACE_LOCATION = "C20R21.le_tile.le_guts.lp0.lut_0";
defparam ii2555.PCK_LOCATION = "C20R21.lp0.lut_0";
defparam ii2555.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2556 (
	. xy ( \ii2556|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2556.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.lut_0";
defparam ii2556.PCK_LOCATION = "C18R22.lp0.lut_0";
defparam ii2556.config_data = 64'b1011000011000000101110111100110010110000110000001011101111001100;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4]|qx_net  ),
	. di ( \ii2491|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .PCK_LOCATION = "C14R9.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_1_In3p_reg[7] .always_en = 1;
LUT6 ii2557 (
	. xy ( \ii2557|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[10]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \ii2555|xy_net  ),
	. f1 ( \carry_13_ADD_10|s_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2557.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.lut_0";
defparam ii2557.PCK_LOCATION = "C18R22.lp0.lut_0";
defparam ii2557.config_data = 64'b1110111100000000111000000000000011101111111011111110000011100000;
LUT6 ii2558 (
	. xy ( \ii2558|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[11]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \ii2555|xy_net  ),
	. f1 ( \carry_13_ADD_11|s_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2558.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.lut_0";
defparam ii2558.PCK_LOCATION = "C18R22.lp0.lut_0";
defparam ii2558.config_data = 64'b1110111100000000111000000000000011101111111011111110000011100000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[13]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[13] .always_en = 1;
LUT6 ii2559 (
	. xy ( \ii2559|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_1|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2559.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2559.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2559.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
LUT6 ii2560 (
	. xy ( \ii2560|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_2|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2560.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2560.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2560.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1]|qx_net  ),
	. di ( \ii2330|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[1] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. di ( \ii2633|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .PCK_LOCATION = "C10R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14] .always_en = 1;
LUT6 ii2561 (
	. xy ( \ii2561|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_3|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2561.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2561.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2561.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_7__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .PCK_LOCATION = "C16R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[0] .always_en = 1;
LUT6 ii2562 (
	. xy ( \ii2562|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_4|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2562.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2562.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2562.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[5] .always_en = 1;
LUT6 ii2563 (
	. xy ( \ii2563|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[5]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_5|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2563.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2563.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2563.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
REG glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload_valid_last_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.PCK_LOCATION = "C4R7.lp0.reg0";
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_rx_payload_valid_last_d_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[18]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .PLACE_LOCATION = "C20R20.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .PCK_LOCATION = "C20R20.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[4] .always_en = 1;
LUT6 ii2564 (
	. xy ( \ii2564|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[6]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_6|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2564.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2564.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2564.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[1]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
LUT6 ii2565 (
	. xy ( \ii2565|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[7]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \carry_13_ADD_7|s_net  ),
	. f1 ( \ii2555|xy_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2565.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2565.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2565.config_data = 64'b1111101100000000110010000000000011111011111110111100100011001000;
REG mcu_arbiter_u_emif2apb_memwr_s_reg (
	. qx ( \mcu_arbiter_u_emif2apb_memwr_s_reg|qx_net  ),
	. di ( \ii3366|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.latch_mode = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.init = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.PLACE_LOCATION = "C4R16.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.sr_inv = 1;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.sync_mode = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.no_sr = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.sr_value = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.PCK_LOCATION = "C4R16.lp0.reg0";
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.clk_inv = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.en_inv = 0;
defparam mcu_arbiter_u_emif2apb_memwr_s_reg.always_en = 1;
LUT6 ii2566 (
	. xy ( \ii2566|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[8]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \ii2555|xy_net  ),
	. f1 ( \carry_13_ADD_8|s_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2566.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.lut_0";
defparam ii2566.PCK_LOCATION = "C18R22.lp0.lut_0";
defparam ii2566.config_data = 64'b1110111100000000111000000000000011101111111011111110000011100000;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5]|qx_net  ),
	. di ( \ii2492|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[5] .always_en = 1;
LUT6 ii2567 (
	. xy ( \ii2567|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t21_out1_reg[9]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f2 ( \ii2555|xy_net  ),
	. f1 ( \carry_13_ADD_9|s_net  ),
	. f0 ( \carry_13_ADD_12|s_net  )
);
defparam ii2567.PLACE_LOCATION = "C18R22.le_tile.le_guts.lp0.lut_0";
defparam ii2567.PCK_LOCATION = "C18R22.lp0.lut_0";
defparam ii2567.config_data = 64'b1110111100000000111000000000000011101111111011111110000011100000;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0]|qx_net  ),
	. di ( \ii2865|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[0] .always_en = 1;
LUT6 ii2568 (
	. xy ( \ii2568|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t24_out1_reg[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2568.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2568.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2568.config_data = 64'b1000110010101111100011001010111110001100101011111000110010101111;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[14]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[14] .always_en = 1;
LUT6 ii2569 (
	. xy ( \ii2569|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_1|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2569.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2569.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2569.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
LUT6 ii2570 (
	. xy ( \ii2570|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_2|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2570.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2570.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2570.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[24]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf.PLACE_LOCATION = "C16R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf.PCK_LOCATION = "C16R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2]|qx_net  ),
	. di ( \ii2331|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[2] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. di ( \ii2637|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .PLACE_LOCATION = "C14R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .PCK_LOCATION = "C14R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15] .always_en = 1;
LUT6 ii2571 (
	. xy ( \ii2571|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_3|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2571.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2571.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2571.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_7__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[1] .always_en = 1;
LUT6 ii2572 (
	. xy ( \ii2572|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_4|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2572.PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.lut_0";
defparam ii2572.PCK_LOCATION = "C20R18.lp0.lut_0";
defparam ii2572.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[6] .always_en = 1;
LUT6 ii2573 (
	. xy ( \ii2573|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_5|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2573.PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.lut_0";
defparam ii2573.PCK_LOCATION = "C18R17.lp0.lut_0";
defparam ii2573.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_4_In1p_reg[5] .always_en = 1;
LUT6 ii2574 (
	. xy ( \ii2574|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_6|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2574.PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.lut_0";
defparam ii2574.PCK_LOCATION = "C20R17.lp0.lut_0";
defparam ii2574.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
LUT6 ii2575 (
	. xy ( \ii2575|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_7|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2575.PLACE_LOCATION = "C20R17.le_tile.le_guts.lp0.lut_0";
defparam ii2575.PCK_LOCATION = "C20R17.lp0.lut_0";
defparam ii2575.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
LUT6 ii2576 (
	. xy ( \ii2576|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_8|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2576.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2576.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2576.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6]|qx_net  ),
	. di ( \ii2493|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[6] .always_en = 1;
LUT6 ii2577 (
	. xy ( \ii2577|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_reg|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t16_out1_reg|qx_net  ),
	. f1 ( \carry_11_ADD_9|s_net  ),
	. f0 ( \carry_11_ADD_10|s_net  )
);
defparam ii2577.PLACE_LOCATION = "C18R18.le_tile.le_guts.lp0.lut_0";
defparam ii2577.PCK_LOCATION = "C18R18.lp0.lut_0";
defparam ii2577.config_data = 64'b1110000011101110111000001110111011100000111011101110000011101110;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1]|qx_net  ),
	. di ( \ii2887|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[1] .always_en = 1;
LUT6 ii2578 (
	. xy ( \ii2578|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2578.PLACE_LOCATION = "C6R15.le_tile.le_guts.lp0.lut_0";
defparam ii2578.PCK_LOCATION = "C6R15.lp0.lut_0";
defparam ii2578.config_data = 64'b1011111001111101000000000000000001000001100000100000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u0_hardfifo_u_inst|dout[15]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[15] .always_en = 1;
LUT6 ii2579 (
	. xy ( \ii2579|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2579.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam ii2579.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam ii2579.config_data = 64'b1110111011110101101011110111011100010001000010100101000010001000;
LUT6 ii2580 (
	. xy ( \ii2580|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]|qx_net  ),
	. f0 ( \ii2579|xy_net  )
);
defparam ii2580.PLACE_LOCATION = "C8R18.le_tile.le_guts.lp0.lut_0";
defparam ii2580.PCK_LOCATION = "C8R18.lp0.lut_0";
defparam ii2580.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3]|qx_net  ),
	. di ( \ii2332|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[3] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. di ( \ii2641|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .PLACE_LOCATION = "C14R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .PCK_LOCATION = "C14R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16] .always_en = 1;
LUT6 ii2581 (
	. xy ( \ii2581|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[1]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[0]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2581.PLACE_LOCATION = "C8R15.le_tile.le_guts.lp0.lut_0";
defparam ii2581.PCK_LOCATION = "C8R15.lp0.lut_0";
defparam ii2581.config_data = 64'b0101000110001010010100001000100001000000100000000000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_7__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[2] .always_en = 1;
LUT6 ii2582 (
	. xy ( \ii2582|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2582.PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.lut_0";
defparam ii2582.PCK_LOCATION = "C14R11.lp0.lut_0";
defparam ii2582.config_data = 64'b1000100010001000100010001000100010001000100010001000100010001000;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .PLACE_LOCATION = "C20R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .PCK_LOCATION = "C20R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[7] .always_en = 1;
LUT6 ii2583 (
	. xy ( \ii2583|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t41_out1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t39_reg_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2581|xy_net  )
);
defparam ii2583.PLACE_LOCATION = "C8R17.le_tile.le_guts.lp0.lut_0";
defparam ii2583.PCK_LOCATION = "C8R17.lp0.lut_0";
defparam ii2583.config_data = 64'b1001010101010101000000000000000001101010101010100000000000000000;
LUT6 ii2584 (
	. xy ( \ii2584|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[0]_net  )
);
defparam ii2584.PLACE_LOCATION = "C20R28.le_tile.le_guts.lp0.lut_0";
defparam ii2584.PCK_LOCATION = "C20R28.lp0.lut_0";
defparam ii2584.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG mcu_arbiter_u_psram_memack_reg (
	. qx ( \mcu_arbiter_u_psram_memack_reg|qx_net  ),
	. di ( \ii3369|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_u_psram_memack_reg.latch_mode = 0;
defparam mcu_arbiter_u_psram_memack_reg.init = 0;
defparam mcu_arbiter_u_psram_memack_reg.PLACE_LOCATION = "C4R18.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_u_psram_memack_reg.sr_inv = 1;
defparam mcu_arbiter_u_psram_memack_reg.sync_mode = 0;
defparam mcu_arbiter_u_psram_memack_reg.no_sr = 0;
defparam mcu_arbiter_u_psram_memack_reg.sr_value = 0;
defparam mcu_arbiter_u_psram_memack_reg.PCK_LOCATION = "C4R18.lp0.reg0";
defparam mcu_arbiter_u_psram_memack_reg.clk_inv = 0;
defparam mcu_arbiter_u_psram_memack_reg.en_inv = 0;
defparam mcu_arbiter_u_psram_memack_reg.always_en = 1;
LUT6 ii2585 (
	. xy ( \ii2585|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[10]_net  )
);
defparam ii2585.PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.lut_0";
defparam ii2585.PCK_LOCATION = "C20R25.lp0.lut_0";
defparam ii2585.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2586 (
	. xy ( \ii2586|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[11]_net  )
);
defparam ii2586.PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.lut_0";
defparam ii2586.PCK_LOCATION = "C20R25.lp0.lut_0";
defparam ii2586.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7]|qx_net  ),
	. di ( \ii2494|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .PCK_LOCATION = "C20R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_5_reg[7] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10]|qx_net  ),
	. di ( \ii2867|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[10] .always_en = 1;
LUT6 ii2587 (
	. xy ( \ii2587|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[12]_net  )
);
defparam ii2587.PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.lut_0";
defparam ii2587.PCK_LOCATION = "C20R25.lp0.lut_0";
defparam ii2587.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
ADD1_A carry_12_0__ADD_10 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[10]|qx_net  ),
	. ci ( \carry_12_0__ADD_9|co_net  ),
	. co ( \carry_12_0__ADD_10|co_net  ),
	. s ( \carry_12_0__ADD_10|s_net  )
);
defparam carry_12_0__ADD_10.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_10.a_inv = "false";
defparam carry_12_0__ADD_10.PCK_LOCATION = "C8R5.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2]|qx_net  ),
	. di ( \ii2909|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[2] .always_en = 1;
LUT6 ii2588 (
	. xy ( \ii2588|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[13]_net  )
);
defparam ii2588.PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.lut_0";
defparam ii2588.PCK_LOCATION = "C20R25.lp0.lut_0";
defparam ii2588.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[16] .always_en = 1;
ADD1_A carry_12_0__ADD_11 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[11]|qx_net  ),
	. ci ( \carry_12_0__ADD_10|co_net  ),
	. co ( ),
	. s ( \carry_12_0__ADD_11|s_net  )
);
defparam carry_12_0__ADD_11.PLACE_LOCATION = "C8R5.le_tile.le_guts.lp0.add2.add0";
defparam carry_12_0__ADD_11.a_inv = "false";
defparam carry_12_0__ADD_11.PCK_LOCATION = "C8R5.lp0.add2.add0";
LUT6 ii2589 (
	. xy ( \ii2589|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[14]_net  )
);
defparam ii2589.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2589.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2589.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2590 (
	. xy ( \ii2590|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[15]_net  )
);
defparam ii2590.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2590.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2590.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2600 (
	. xy ( \ii2600|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[2]_net  )
);
defparam ii2600.PLACE_LOCATION = "C20R27.le_tile.le_guts.lp0.lut_0";
defparam ii2600.PCK_LOCATION = "C20R27.lp0.lut_0";
defparam ii2600.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4]|qx_net  ),
	. di ( \ii2333|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[4] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. di ( \ii2646|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17] .always_en = 1;
LUT6 ii2591 (
	. xy ( \ii2591|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[16]_net  )
);
defparam ii2591.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2591.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2591.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2601 (
	. xy ( \ii2601|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[3]_net  )
);
defparam ii2601.PLACE_LOCATION = "C20R28.le_tile.le_guts.lp0.lut_0";
defparam ii2601.PCK_LOCATION = "C20R28.lp0.lut_0";
defparam ii2601.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3]|qx_net  ),
	. di ( \carry_9_7__ADD_3|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .PLACE_LOCATION = "C18R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .PCK_LOCATION = "C18R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[3] .always_en = 1;
LUT6 ii2592 (
	. xy ( \ii2592|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[17]_net  )
);
defparam ii2592.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2592.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2592.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2602 (
	. xy ( \ii2602|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[4]_net  )
);
defparam ii2602.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2602.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2602.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .PLACE_LOCATION = "C16R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .PCK_LOCATION = "C16R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[8] .always_en = 1;
LUT6 ii2593 (
	. xy ( \ii2593|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[18]_net  )
);
defparam ii2593.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2593.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2593.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2603 (
	. xy ( \ii2603|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[5]_net  )
);
defparam ii2603.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2603.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2603.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2594 (
	. xy ( \ii2594|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[19]_net  )
);
defparam ii2594.PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.lut_0";
defparam ii2594.PCK_LOCATION = "C16R26.lp0.lut_0";
defparam ii2594.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2604 (
	. xy ( \ii2604|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[6]_net  )
);
defparam ii2604.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2604.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2604.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2595 (
	. xy ( \ii2595|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[1]_net  )
);
defparam ii2595.PLACE_LOCATION = "C20R28.le_tile.le_guts.lp0.lut_0";
defparam ii2595.PCK_LOCATION = "C20R28.lp0.lut_0";
defparam ii2595.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2605 (
	. xy ( \ii2605|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[7]_net  )
);
defparam ii2605.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2605.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2605.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf (
	. xy ( \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( ),
	. f0 ( \mcu_arbiter_u_emif2apb_write_data_temp_reg[14]|qx_net  )
);
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf.PLACE_LOCATION = "C14R14.le_tile.le_guts.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf.PCK_LOCATION = "C14R14.lp0.lut_0";
defparam mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf.config_data = 64'b1010101010101010101010101010101010101010101010101010101010101010;
REG \mcu_arbiter_u_psram_dsel_reg[0]  (
	. qx ( \mcu_arbiter_u_psram_dsel_reg[0]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memaddr_comb[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_psram_dsel_reg[0] .latch_mode = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .init = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_psram_dsel_reg[0] .sr_inv = 1;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .sync_mode = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .no_sr = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .sr_value = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \mcu_arbiter_u_psram_dsel_reg[0] .clk_inv = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .en_inv = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[0] .always_en = 1;
LUT6 ii2596 (
	. xy ( \ii2596|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[20]_net  )
);
defparam ii2596.PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.lut_0";
defparam ii2596.PCK_LOCATION = "C16R26.lp0.lut_0";
defparam ii2596.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2606 (
	. xy ( \ii2606|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[8]_net  )
);
defparam ii2606.PLACE_LOCATION = "C18R25.le_tile.le_guts.lp0.lut_0";
defparam ii2606.PCK_LOCATION = "C18R25.lp0.lut_0";
defparam ii2606.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11]|qx_net  ),
	. di ( \ii2869|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[11] .always_en = 1;
LUT6 ii2597 (
	. xy ( \ii2597|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[21]_net  )
);
defparam ii2597.PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.lut_0";
defparam ii2597.PCK_LOCATION = "C16R26.lp0.lut_0";
defparam ii2597.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2607 (
	. xy ( \ii2607|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[9]_net  )
);
defparam ii2607.PLACE_LOCATION = "C20R25.le_tile.le_guts.lp0.lut_0";
defparam ii2607.PCK_LOCATION = "C20R25.lp0.lut_0";
defparam ii2607.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3]|qx_net  ),
	. di ( \ii2915|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[3] .always_en = 1;
LUT6 ii2598 (
	. xy ( \ii2598|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[22]_net  )
);
defparam ii2598.PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.lut_0";
defparam ii2598.PCK_LOCATION = "C16R26.lp0.lut_0";
defparam ii2598.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2608 (
	. xy ( \ii2608|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_reg|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t13_out1_reg|qx_net  ),
	. f0 ( \ii2555|xy_net  )
);
defparam ii2608.PLACE_LOCATION = "C20R22.le_tile.le_guts.lp0.lut_0";
defparam ii2608.PCK_LOCATION = "C20R22.lp0.lut_0";
defparam ii2608.config_data = 64'b1011101010111010101110101011101010111010101110101011101010111010;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[17] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[0] .always_en = 1;
LUT6 ii2599 (
	. xy ( \ii2599|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t50_out1_reg|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_u_emb1_xx2_u_spram|datao[23]_net  )
);
defparam ii2599.PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.lut_0";
defparam ii2599.PCK_LOCATION = "C16R26.lp0.lut_0";
defparam ii2599.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
LUT6 ii2609 (
	. xy ( \ii2609|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  )
);
defparam ii2609.PLACE_LOCATION = "C10R10.le_tile.le_guts.lp0.lut_0";
defparam ii2609.PCK_LOCATION = "C10R10.lp0.lut_0";
defparam ii2609.config_data = 64'b0001000100010001000100010001000100010001000100010001000100010001;
LUT6 ii2610 (
	. xy ( \ii2610|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[0]|qx_net  )
);
defparam ii2610.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2610.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2610.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
SIO io_rx_decode_vsync_inst (
	. f_id ( )
,
	. clk_en ( ),
	. fclk ( ),
	. od ( {
		/* od [1] (nc) */ nc569 ,
		/* od [0] */ \glue_rx_packet_tx_packet_u_data_process_fifo_writeen_reg|qx_net 
	} ),
	. oen ( ),
	. rstn ( ),
	. setn ( ),
	. PAD ( rx_decode_vsync )
);
defparam io_rx_decode_vsync_inst.DDR_PREG_EN = 0;
defparam io_rx_decode_vsync_inst.FCLK_GATE_EN = 0;
defparam io_rx_decode_vsync_inst.FOEN_SEL = 0;
defparam io_rx_decode_vsync_inst.RSTN_SYNC = 0;
defparam io_rx_decode_vsync_inst.OUT_SEL = 2;
defparam io_rx_decode_vsync_inst.DDR_EN = 0;
defparam io_rx_decode_vsync_inst.NDR = 15;
defparam io_rx_decode_vsync_inst.VPCI_EN = 0;
defparam io_rx_decode_vsync_inst.ID_RSTN_EN = 0;
defparam io_rx_decode_vsync_inst.KEEP = 0;
defparam io_rx_decode_vsync_inst.PDR = 15;
defparam io_rx_decode_vsync_inst.SETN_INV = 0;
defparam io_rx_decode_vsync_inst.SETN_SYNC = 0;
defparam io_rx_decode_vsync_inst.FIN_SEL = 0;
defparam io_rx_decode_vsync_inst.ID_SETN_EN = 0;
defparam io_rx_decode_vsync_inst.DDR_REG_EN = 0;
defparam io_rx_decode_vsync_inst.FOUT_SEL = 0;
defparam io_rx_decode_vsync_inst.OEN_RSTN_EN = 0;
defparam io_rx_decode_vsync_inst.NS_LV = 3;
defparam io_rx_decode_vsync_inst.optional_function = "";
defparam io_rx_decode_vsync_inst.OD_RSTN_EN = 0;
defparam io_rx_decode_vsync_inst.RSTN_INV = 0;
defparam io_rx_decode_vsync_inst.is_clk_io = "false";
defparam io_rx_decode_vsync_inst.PLACE_LOCATION = "C24R17.io_guts.iob_ck.I0.I60.Iioc1";
defparam io_rx_decode_vsync_inst.OEN_SETN_EN = 0;
defparam io_rx_decode_vsync_inst.OEN_SEL = 1;
defparam io_rx_decode_vsync_inst.PCK_LOCATION = "NONE";
defparam io_rx_decode_vsync_inst.OD_SETN_EN = 0;
defparam io_rx_decode_vsync_inst.CLK_INV = 0;
defparam io_rx_decode_vsync_inst.is_signal_monitor_io = 1'b0;
defparam io_rx_decode_vsync_inst.DDR_NREG_EN = 0;
defparam io_rx_decode_vsync_inst.RX_DIG_EN = 0;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5]|qx_net  ),
	. di ( \ii2334|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[5] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. di ( \ii2651|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18] .always_en = 1;
LUT6 ii2611 (
	. xy ( \ii2611|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]|qx_net  ),
	. f1 ( \ii2610|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2611.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2611.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2611.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4]|qx_net  ),
	. di ( \carry_9_7__ADD_4|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[4] .always_en = 1;
LUT6 ii2612 (
	. xy ( \ii2612|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  )
);
defparam ii2612.PLACE_LOCATION = "C14R11.le_tile.le_guts.lp0.lut_0";
defparam ii2612.PCK_LOCATION = "C14R11.lp0.lut_0";
defparam ii2612.config_data = 64'b0010001000100010001000100010001000100010001000100010001000100010;
REG \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t6_out1_reg[9]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .PLACE_LOCATION = "C20R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .PCK_LOCATION = "C20R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[9] .always_en = 1;
LUT6 ii2613 (
	. xy ( \ii2613|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[0]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2611|xy_net  )
);
defparam ii2613.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2613.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2613.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_sync_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_frame_start_d_reg.always_en = 1;
LUT6 ii2614 (
	. xy ( \ii2614|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2614.PLACE_LOCATION = "C10R8.le_tile.le_guts.lp0.lut_0";
defparam ii2614.PCK_LOCATION = "C10R8.lp0.lut_0";
defparam ii2614.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
MIPI_TOP mipi_inst_u_mipi1 (
	. CN ( )
,
	. CM ( )
,
	. CO ( )
,
	. port_sel ( {
		/* port_sel [1] */ \VCC_0_inst|Y_net ,
		/* port_sel [0] */ \GND_0_inst|Y_net 
	} ),
	. enable_raw_dsi_port ( \VCC_0_inst|Y_net  ),
	. enable_dpi_port ( \GND_0_inst|Y_net  ),
	. TxEscClk ( \u_pll_pll_u0|CO1_net  ),
	. RxEscClk ( \u_pll_pll_u0|CO2_net  ),
	. reset_n ( \ii2048|xy_net  ),
	. reset_esc_n ( \ii2048|xy_net  ),
	. clk_periph ( \u_pll_pll_u0|CO0_net  ),
	. RxSyncHS ( ),
	. RxActiveHS ( \mipi_inst_u_mipi1|RxActiveHS_net  ),
	. RxLpdtEsc ( ),
	. periph_dpi_vsync ( ),
	. periph_dpi_hsync ( ),
	. periph_dpi_de ( ),
	. periph_dpi_d ( )
,
	. periph_dpi_sd ( ),
	. periph_dpi_cm ( ),
	. periph_dpi_peripheral_output_dropped ( ),
	. periph_rx_cmd ( {
		/* periph_rx_cmd [23] (nc) */ nc570 ,
		/* periph_rx_cmd [22] (nc) */ nc571 ,
		/* periph_rx_cmd [21] (nc) */ nc572 ,
		/* periph_rx_cmd [20] (nc) */ nc573 ,
		/* periph_rx_cmd [19] (nc) */ nc574 ,
		/* periph_rx_cmd [18] (nc) */ nc575 ,
		/* periph_rx_cmd [17] (nc) */ nc576 ,
		/* periph_rx_cmd [16] (nc) */ nc577 ,
		/* periph_rx_cmd [15] */ \mipi_inst_u_mipi1|periph_rx_cmd[15]_net ,
		/* periph_rx_cmd [14] */ \mipi_inst_u_mipi1|periph_rx_cmd[14]_net ,
		/* periph_rx_cmd [13] */ \mipi_inst_u_mipi1|periph_rx_cmd[13]_net ,
		/* periph_rx_cmd [12] */ \mipi_inst_u_mipi1|periph_rx_cmd[12]_net ,
		/* periph_rx_cmd [11] */ \mipi_inst_u_mipi1|periph_rx_cmd[11]_net ,
		/* periph_rx_cmd [10] */ \mipi_inst_u_mipi1|periph_rx_cmd[10]_net ,
		/* periph_rx_cmd [9] */ \mipi_inst_u_mipi1|periph_rx_cmd[9]_net ,
		/* periph_rx_cmd [8] */ \mipi_inst_u_mipi1|periph_rx_cmd[8]_net ,
		/* periph_rx_cmd [7] (nc) */ nc578 ,
		/* periph_rx_cmd [6] (nc) */ nc579 ,
		/* periph_rx_cmd [5] */ \mipi_inst_u_mipi1|periph_rx_cmd[5]_net ,
		/* periph_rx_cmd [4] */ \mipi_inst_u_mipi1|periph_rx_cmd[4]_net ,
		/* periph_rx_cmd [3] */ \mipi_inst_u_mipi1|periph_rx_cmd[3]_net ,
		/* periph_rx_cmd [2] */ \mipi_inst_u_mipi1|periph_rx_cmd[2]_net ,
		/* periph_rx_cmd [1] */ \mipi_inst_u_mipi1|periph_rx_cmd[1]_net ,
		/* periph_rx_cmd [0] */ \mipi_inst_u_mipi1|periph_rx_cmd[0]_net 
	} ),
	. periph_rx_cmd_valid ( \mipi_inst_u_mipi1|periph_rx_cmd_valid_net  ),
	. periph_rx_payload ( {
		/* periph_rx_payload [31] */ \mipi_inst_u_mipi1|periph_rx_payload[31]_net ,
		/* periph_rx_payload [30] */ \mipi_inst_u_mipi1|periph_rx_payload[30]_net ,
		/* periph_rx_payload [29] */ \mipi_inst_u_mipi1|periph_rx_payload[29]_net ,
		/* periph_rx_payload [28] */ \mipi_inst_u_mipi1|periph_rx_payload[28]_net ,
		/* periph_rx_payload [27] */ \mipi_inst_u_mipi1|periph_rx_payload[27]_net ,
		/* periph_rx_payload [26] */ \mipi_inst_u_mipi1|periph_rx_payload[26]_net ,
		/* periph_rx_payload [25] */ \mipi_inst_u_mipi1|periph_rx_payload[25]_net ,
		/* periph_rx_payload [24] */ \mipi_inst_u_mipi1|periph_rx_payload[24]_net ,
		/* periph_rx_payload [23] */ \mipi_inst_u_mipi1|periph_rx_payload[23]_net ,
		/* periph_rx_payload [22] */ \mipi_inst_u_mipi1|periph_rx_payload[22]_net ,
		/* periph_rx_payload [21] */ \mipi_inst_u_mipi1|periph_rx_payload[21]_net ,
		/* periph_rx_payload [20] */ \mipi_inst_u_mipi1|periph_rx_payload[20]_net ,
		/* periph_rx_payload [19] */ \mipi_inst_u_mipi1|periph_rx_payload[19]_net ,
		/* periph_rx_payload [18] */ \mipi_inst_u_mipi1|periph_rx_payload[18]_net ,
		/* periph_rx_payload [17] */ \mipi_inst_u_mipi1|periph_rx_payload[17]_net ,
		/* periph_rx_payload [16] */ \mipi_inst_u_mipi1|periph_rx_payload[16]_net ,
		/* periph_rx_payload [15] */ \mipi_inst_u_mipi1|periph_rx_payload[15]_net ,
		/* periph_rx_payload [14] */ \mipi_inst_u_mipi1|periph_rx_payload[14]_net ,
		/* periph_rx_payload [13] */ \mipi_inst_u_mipi1|periph_rx_payload[13]_net ,
		/* periph_rx_payload [12] */ \mipi_inst_u_mipi1|periph_rx_payload[12]_net ,
		/* periph_rx_payload [11] */ \mipi_inst_u_mipi1|periph_rx_payload[11]_net ,
		/* periph_rx_payload [10] */ \mipi_inst_u_mipi1|periph_rx_payload[10]_net ,
		/* periph_rx_payload [9] */ \mipi_inst_u_mipi1|periph_rx_payload[9]_net ,
		/* periph_rx_payload [8] */ \mipi_inst_u_mipi1|periph_rx_payload[8]_net ,
		/* periph_rx_payload [7] */ \mipi_inst_u_mipi1|periph_rx_payload[7]_net ,
		/* periph_rx_payload [6] */ \mipi_inst_u_mipi1|periph_rx_payload[6]_net ,
		/* periph_rx_payload [5] */ \mipi_inst_u_mipi1|periph_rx_payload[5]_net ,
		/* periph_rx_payload [4] */ \mipi_inst_u_mipi1|periph_rx_payload[4]_net ,
		/* periph_rx_payload [3] */ \mipi_inst_u_mipi1|periph_rx_payload[3]_net ,
		/* periph_rx_payload [2] */ \mipi_inst_u_mipi1|periph_rx_payload[2]_net ,
		/* periph_rx_payload [1] */ \mipi_inst_u_mipi1|periph_rx_payload[1]_net ,
		/* periph_rx_payload [0] */ \mipi_inst_u_mipi1|periph_rx_payload[0]_net 
	} ),
	. periph_rx_payload_valid ( \mipi_inst_u_mipi1|periph_rx_payload_valid_net  ),
	. periph_rx_payload_valid_last ( \mipi_inst_u_mipi1|periph_rx_payload_valid_last_net  ),
	. periph_rx_trigger ( )
,
	. periph_rx_trigger_valid ( ),
	. periph_ecc_one_bit_err ( ),
	. periph_ecc_two_bit_err ( ),
	. periph_ecc_one_bit_err_pos ( )
,
	. periph_ecc_err ( ),
	. periph_ecc_err_pos ( )
,
	. periph_crc_err ( ),
	. periph_te_enable ( \GND_0_inst|Y_net  ),
	. periph_te_rdy ( ),
	. periph_te_ack ( ),
	. periph_te_event_in ( \GND_0_inst|Y_net  ),
	. periph_te_fail ( \GND_0_inst|Y_net  ),
	. periph_rx_ulps_active ( )
,
	. periph_rx_ulps_mark_active ( )
,
	. periph_tx_payload ( {
		/* periph_tx_payload [31] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[31]|qx_net ,
		/* periph_tx_payload [30] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[30]|qx_net ,
		/* periph_tx_payload [29] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[29]|qx_net ,
		/* periph_tx_payload [28] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[28]|qx_net ,
		/* periph_tx_payload [27] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[27]|qx_net ,
		/* periph_tx_payload [26] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[26]|qx_net ,
		/* periph_tx_payload [25] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[25]|qx_net ,
		/* periph_tx_payload [24] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[24]|qx_net ,
		/* periph_tx_payload [23] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[23]|qx_net ,
		/* periph_tx_payload [22] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[22]|qx_net ,
		/* periph_tx_payload [21] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[21]|qx_net ,
		/* periph_tx_payload [20] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[20]|qx_net ,
		/* periph_tx_payload [19] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[19]|qx_net ,
		/* periph_tx_payload [18] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[18]|qx_net ,
		/* periph_tx_payload [17] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[17]|qx_net ,
		/* periph_tx_payload [16] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[16]|qx_net ,
		/* periph_tx_payload [15] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[15]|qx_net ,
		/* periph_tx_payload [14] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[14]|qx_net ,
		/* periph_tx_payload [13] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[13]|qx_net ,
		/* periph_tx_payload [12] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[12]|qx_net ,
		/* periph_tx_payload [11] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[11]|qx_net ,
		/* periph_tx_payload [10] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[10]|qx_net ,
		/* periph_tx_payload [9] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[9]|qx_net ,
		/* periph_tx_payload [8] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[8]|qx_net ,
		/* periph_tx_payload [7] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[7]|qx_net ,
		/* periph_tx_payload [6] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[6]|qx_net ,
		/* periph_tx_payload [5] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[5]|qx_net ,
		/* periph_tx_payload [4] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[4]|qx_net ,
		/* periph_tx_payload [3] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[3]|qx_net ,
		/* periph_tx_payload [2] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[2]|qx_net ,
		/* periph_tx_payload [1] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[1]|qx_net ,
		/* periph_tx_payload [0] */ \uut_dataReadBack_mipi_periph_tx_payload_reg[0]|qx_net 
	} ),
	. periph_tx_payload_en ( ),
	. periph_tx_payload_en_last ( ),
	. periph_tx_cmd_vc ( {
		/* periph_tx_cmd_vc [1] */ \GND_0_inst|Y_net ,
		/* periph_tx_cmd_vc [0] */ \GND_0_inst|Y_net 
	} ),
	. periph_tx_cmd_data_type ( {
		/* periph_tx_cmd_data_type [5] */ \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[5]|qx_net ,
		/* periph_tx_cmd_data_type [4] */ \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[4]|qx_net ,
		/* periph_tx_cmd_data_type [3] */ \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[3]|qx_net ,
		/* periph_tx_cmd_data_type [2] */ \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[2]|qx_net ,
		/* periph_tx_cmd_data_type [1] */ \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[1]|qx_net ,
		/* periph_tx_cmd_data_type [0] */ \uut_dataReadBack_mipi_periph_tx_cmd_data_type_reg[0]|qx_net 
	} ),
	. periph_tx_cmd_byte_count ( {
		/* periph_tx_cmd_byte_count [15] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[15]|qx_net ,
		/* periph_tx_cmd_byte_count [14] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[14]|qx_net ,
		/* periph_tx_cmd_byte_count [13] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[13]|qx_net ,
		/* periph_tx_cmd_byte_count [12] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[12]|qx_net ,
		/* periph_tx_cmd_byte_count [11] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[11]|qx_net ,
		/* periph_tx_cmd_byte_count [10] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[10]|qx_net ,
		/* periph_tx_cmd_byte_count [9] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[9]|qx_net ,
		/* periph_tx_cmd_byte_count [8] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[8]|qx_net ,
		/* periph_tx_cmd_byte_count [7] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[7]|qx_net ,
		/* periph_tx_cmd_byte_count [6] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[6]|qx_net ,
		/* periph_tx_cmd_byte_count [5] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[5]|qx_net ,
		/* periph_tx_cmd_byte_count [4] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[4]|qx_net ,
		/* periph_tx_cmd_byte_count [3] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[3]|qx_net ,
		/* periph_tx_cmd_byte_count [2] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[2]|qx_net ,
		/* periph_tx_cmd_byte_count [1] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[1]|qx_net ,
		/* periph_tx_cmd_byte_count [0] */ \uut_dataReadBack_mipi_periph_tx_cmd_byte_count_reg[0]|qx_net 
	} ),
	. periph_tx_cmd_req ( \uut_dataReadBack_mipi_periph_tx_cmd_req_reg|qx_net  ),
	. periph_tx_cmd_ack ( \mipi_inst_u_mipi1|periph_tx_cmd_ack_net  ),
	. periph_tx_timeout_error ( ),
	. periph_trigger_req ( \GND_0_inst|Y_net  ),
	. periph_trigger_ack ( ),
	. periph_trigger_send ( {
		/* periph_trigger_send [1] */ \GND_0_inst|Y_net ,
		/* periph_trigger_send [0] */ \GND_0_inst|Y_net 
	} ),
	. periph_dphy_direction ( \mipi_inst_u_mipi1|periph_dphy_direction_net  ),
	. hs_rx_timeout ( ),
	. lp_tx_timeout ( ),
	. periph_bta_timeout ( ),
	. dpi_pclk ( ),
	. reset_dpi_n ( ),
	. host_dpi_vsync ( ),
	. host_dpi_hsync ( ),
	. host_dpi_de ( ),
	. host_dpi_d ( )
,
	. host_dpi_sd ( ),
	. host_dpi_cm ( ),
	. dpi_host_underrun_err ( ),
	. host_tx_cmd_vc ( )
,
	. host_tx_cmd_data_type ( )
,
	. host_tx_cmd_byte_count ( )
,
	. host_tx_cmd_ack ( ),
	. host_tx_cmd_req ( ),
	. host_tx_payload ( )
,
	. host_tx_payload_en ( ),
	. host_tx_payload_en_last ( ),
	. host_tx_hs_mode ( ),
	. host_tx_active ( ),
	. host_tx_ulps_enable ( )
,
	. host_tx_ulps_active ( )
,
	. host_dphy_turnaround ( ),
	. host_dphy_direction ( ),
	. host_trigger_req ( ),
	. host_trigger_send ( )
,
	. host_trigger_ack ( ),
	. host_rx_payload ( )
,
	. host_rx_payload_valid ( ),
	. host_rx_payload_valid_last ( ),
	. host_rx_cmd_valid ( ),
	. host_rx_cmd_vc ( )
,
	. host_rx_cmd_data_type ( )
,
	. host_rx_cmd_byte_count ( )
,
	. host_ecc_one_bit_err ( ),
	. host_ecc_two_bit_err ( ),
	. host_ecc_one_bit_err_pos ( )
,
	. host_ecc_err ( ),
	. host_ecc_err_pos ( )
,
	. host_crc_err ( ),
	. host_hs_tx_timeout ( ),
	. host_lp_rx_timeout ( ),
	. host_bta_timeout ( ),
	. pclk_reset_n ( \ii1982|xy_net  ),
	. pclk ( \u_pll_pll_u0|CO3_net  ),
	. paddr ( {
		/* paddr [17] */ \GND_0_inst|Y_net ,
		/* paddr [16] */ \GND_0_inst|Y_net ,
		/* paddr [15] */ \GND_0_inst|Y_net ,
		/* paddr [14] */ \GND_0_inst|Y_net ,
		/* paddr [13] */ \GND_0_inst|Y_net ,
		/* paddr [12] */ \GND_0_inst|Y_net ,
		/* paddr [11] */ \GND_0_inst|Y_net ,
		/* paddr [10] */ \GND_0_inst|Y_net ,
		/* paddr [9] */ \u_8051_u_h6_8051|memaddr_comb[9]_net ,
		/* paddr [8] */ \u_8051_u_h6_8051|memaddr_comb[8]_net ,
		/* paddr [7] */ \u_8051_u_h6_8051|memaddr_comb[7]_net ,
		/* paddr [6] */ \u_8051_u_h6_8051|memaddr_comb[6]_net ,
		/* paddr [5] */ \u_8051_u_h6_8051|memaddr_comb[5]_net ,
		/* paddr [4] */ \u_8051_u_h6_8051|memaddr_comb[4]_net ,
		/* paddr [3] */ \u_8051_u_h6_8051|memaddr_comb[3]_net ,
		/* paddr [2] */ \u_8051_u_h6_8051|memaddr_comb[2]_net ,
		/* paddr [1] */ \GND_0_inst|Y_net ,
		/* paddr [0] */ \GND_0_inst|Y_net 
	} ),
	. pwrite ( \mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf|xy_net  ),
	. psel ( \ii2051|xy_net  ),
	. penable ( \ii2050|xy_net  ),
	. pwdata ( {
		/* pwdata [31] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf|xy_net ,
		/* pwdata [30] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf|xy_net ,
		/* pwdata [29] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf|xy_net ,
		/* pwdata [28] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf|xy_net ,
		/* pwdata [27] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf|xy_net ,
		/* pwdata [26] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf|xy_net ,
		/* pwdata [25] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf|xy_net ,
		/* pwdata [24] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf|xy_net ,
		/* pwdata [23] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf|xy_net ,
		/* pwdata [22] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf|xy_net ,
		/* pwdata [21] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf|xy_net ,
		/* pwdata [20] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf|xy_net ,
		/* pwdata [19] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf|xy_net ,
		/* pwdata [18] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf|xy_net ,
		/* pwdata [17] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf|xy_net ,
		/* pwdata [16] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf|xy_net ,
		/* pwdata [15] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf|xy_net ,
		/* pwdata [14] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf|xy_net ,
		/* pwdata [13] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf|xy_net ,
		/* pwdata [12] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf|xy_net ,
		/* pwdata [11] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf|xy_net ,
		/* pwdata [10] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf|xy_net ,
		/* pwdata [9] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf|xy_net ,
		/* pwdata [8] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf|xy_net ,
		/* pwdata [7] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf|xy_net ,
		/* pwdata [6] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf|xy_net ,
		/* pwdata [5] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf|xy_net ,
		/* pwdata [4] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf|xy_net ,
		/* pwdata [3] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf|xy_net ,
		/* pwdata [2] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf|xy_net ,
		/* pwdata [1] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf|xy_net ,
		/* pwdata [0] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf|xy_net 
	} ),
	. prdata ( {
		/* prdata [31] */ \mipi_inst_u_mipi1|prdata[31]_net ,
		/* prdata [30] */ \mipi_inst_u_mipi1|prdata[30]_net ,
		/* prdata [29] */ \mipi_inst_u_mipi1|prdata[29]_net ,
		/* prdata [28] */ \mipi_inst_u_mipi1|prdata[28]_net ,
		/* prdata [27] */ \mipi_inst_u_mipi1|prdata[27]_net ,
		/* prdata [26] */ \mipi_inst_u_mipi1|prdata[26]_net ,
		/* prdata [25] */ \mipi_inst_u_mipi1|prdata[25]_net ,
		/* prdata [24] */ \mipi_inst_u_mipi1|prdata[24]_net ,
		/* prdata [23] */ \mipi_inst_u_mipi1|prdata[23]_net ,
		/* prdata [22] */ \mipi_inst_u_mipi1|prdata[22]_net ,
		/* prdata [21] */ \mipi_inst_u_mipi1|prdata[21]_net ,
		/* prdata [20] */ \mipi_inst_u_mipi1|prdata[20]_net ,
		/* prdata [19] */ \mipi_inst_u_mipi1|prdata[19]_net ,
		/* prdata [18] */ \mipi_inst_u_mipi1|prdata[18]_net ,
		/* prdata [17] */ \mipi_inst_u_mipi1|prdata[17]_net ,
		/* prdata [16] */ \mipi_inst_u_mipi1|prdata[16]_net ,
		/* prdata [15] */ \mipi_inst_u_mipi1|prdata[15]_net ,
		/* prdata [14] */ \mipi_inst_u_mipi1|prdata[14]_net ,
		/* prdata [13] */ \mipi_inst_u_mipi1|prdata[13]_net ,
		/* prdata [12] */ \mipi_inst_u_mipi1|prdata[12]_net ,
		/* prdata [11] */ \mipi_inst_u_mipi1|prdata[11]_net ,
		/* prdata [10] */ \mipi_inst_u_mipi1|prdata[10]_net ,
		/* prdata [9] */ \mipi_inst_u_mipi1|prdata[9]_net ,
		/* prdata [8] */ \mipi_inst_u_mipi1|prdata[8]_net ,
		/* prdata [7] */ \mipi_inst_u_mipi1|prdata[7]_net ,
		/* prdata [6] */ \mipi_inst_u_mipi1|prdata[6]_net ,
		/* prdata [5] */ \mipi_inst_u_mipi1|prdata[5]_net ,
		/* prdata [4] */ \mipi_inst_u_mipi1|prdata[4]_net ,
		/* prdata [3] */ \mipi_inst_u_mipi1|prdata[3]_net ,
		/* prdata [2] */ \mipi_inst_u_mipi1|prdata[2]_net ,
		/* prdata [1] */ \mipi_inst_u_mipi1|prdata[1]_net ,
		/* prdata [0] */ \mipi_inst_u_mipi1|prdata[0]_net 
	} ),
	. pready ( \mipi_inst_u_mipi1|pready_net  ),
	. clk ( ),
	. RxByteClkHS ( ),
	. CLKP ( ),
	. CLKN ( ),
	. DATAN0 ( ),
	. DATAP0 ( ),
	. DATAN1 ( ),
	. DATAP1 ( ),
	. DATAN2 ( ),
	. DATAP2 ( ),
	. DATAN3 ( ),
	. DATAP3 ( ),
	. LOCK ( ),
	. BITCLK ( \mipi_inst_u_mipi_pll|CLKOUT1_net  ),
	. PD_DPHY ( \ii2049|xy_net  ),
	. ENP_DESER ( \GND_0_inst|Y_net  ),
	. TEST_ENBL ( {
		/* TEST_ENBL [5] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [4] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [3] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [2] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [1] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [0] */ \GND_0_inst|Y_net 
	} ),
	. TEST_PATTERN ( )
,
	. D0_LB_PASS ( )
,
	. D1_LB_PASS ( )
,
	. D2_LB_PASS ( )
,
	. D3_LB_PASS ( )
,
	. D0_LB_ERR_CNT ( )
,
	. D1_LB_ERR_CNT ( )
,
	. D2_LB_ERR_CNT ( )
,
	. D3_LB_ERR_CNT ( )
,
	. D0_LB_BYTE_CNT ( )
,
	. D1_LB_BYTE_CNT ( )
,
	. D2_LB_BYTE_CNT ( )
,
	. D3_LB_BYTE_CNT ( )
,
	. D0_LB_ACTIVE ( )
,
	. D1_LB_ACTIVE ( )
,
	. D2_LB_ACTIVE ( )
,
	. D3_LB_ACTIVE ( )
,
	. D0_LB_VALID ( )
,
	. D1_LB_VALID ( )
,
	. D2_LB_VALID ( )
,
	. D3_LB_VALID ( )
,
	. CLK_LB_ACTIVE ( ),
	. DC_TEST_OUT ( )
,
	. AUTO_PD_EN ( \GND_0_inst|Y_net  ),
	. ext_TxRequestHS_lnclk ( ),
	. Stopstate_lnclk ( ),
	. ext_TxUlpsClk_lnclk ( ),
	. ext_TxUlpsExit_lnclk ( ),
	. UlpsActiveNot_lnclk ( ),
	. RxUlpsClkNot ( ),
	. RxClkActiveHS ( ),
	. ext_Enable_lnclk ( ),
	. ext_TxDataHS_ln0 ( )
,
	. ext_TxRequestHS_ln0 ( ),
	. TxReadyHS_ln0 ( ),
	. ext_Enable_ln0 ( ),
	. ext_TxRequestEsc_ln0 ( ),
	. ext_TxUlpsEsc_ln0 ( ),
	. ext_TxLpdtEsc_ln0 ( ),
	. ext_TxUlpsExit_ln0 ( ),
	. TxReadyEsc_ln0 ( ),
	. ext_TxTriggerEsc_ln0 ( )
,
	. ext_TxDataEsc_ln0 ( )
,
	. ext_TxValidEsc_ln0 ( ),
	. ext_ForceTxStopmode_ln0 ( ),
	. ext_TurnRequest_ln0 ( ),
	. ext_TurnDisable_ln0 ( ),
	. ext_ForceRxmode_ln0 ( ),
	. RxClkEsc_ln0 ( ),
	. RxLpdtEsc_ln0 ( ),
	. RxUlpsEsc_ln0 ( ),
	. RxTriggerEsc_ln0 ( )
,
	. RxDataEsc_ln0 ( )
,
	. RxValidEsc_ln0 ( ),
	. Direction_ln0 ( ),
	. Stopstate_ln0 ( ),
	. UlpsActiveNot_ln0 ( ),
	. ErrSotHS_ln0 ( ),
	. ErrSotSyncHS_ln0 ( ),
	. ErrEsc_ln0 ( ),
	. ErrSyncEsc_ln0 ( ),
	. ErrControl_ln0 ( ),
	. ErrContentionLp0_ln0 ( ),
	. ErrContentionLp1_ln0 ( ),
	. RxDataHS_ln0 ( )
,
	. RxValidHS_ln0 ( ),
	. RxActiveHS_ln0 ( ),
	. RxSyncHS_ln0 ( ),
	. ext_TxDataHS_ln1 ( )
,
	. ext_TxRequestHS_ln1 ( ),
	. TxReadyHS_ln1 ( ),
	. ext_Enable_ln1 ( ),
	. ext_TxRequestEsc_ln1 ( ),
	. ext_TxUlpsEsc_ln1 ( ),
	. ext_TxLpdtEsc_ln1 ( ),
	. ext_TxUlpsExit_ln1 ( ),
	. TxReadyEsc_ln1 ( ),
	. ext_TxTriggerEsc_ln1 ( )
,
	. ext_TxDataEsc_ln1 ( )
,
	. ext_TxValidEsc_ln1 ( ),
	. ext_ForceTxStopmode_ln1 ( ),
	. ext_TurnRequest_ln1 ( ),
	. ext_TurnDisable_ln1 ( ),
	. ext_ForceRxmode_ln1 ( ),
	. RxClkEsc_ln1 ( ),
	. RxLpdtEsc_ln1 ( ),
	. RxUlpsEsc_ln1 ( ),
	. RxTriggerEsc_ln1 ( )
,
	. RxDataEsc_ln1 ( )
,
	. RxValidEsc_ln1 ( ),
	. Direction_ln1 ( ),
	. Stopstate_ln1 ( ),
	. UlpsActiveNot_ln1 ( ),
	. ErrSotHS_ln1 ( ),
	. ErrSotSyncHS_ln1 ( ),
	. ErrEsc_ln1 ( ),
	. ErrSyncEsc_ln1 ( ),
	. ErrControl_ln1 ( ),
	. ErrContentionLp0_ln1 ( ),
	. ErrContentionLp1_ln1 ( ),
	. RxDataHS_ln1 ( )
,
	. RxValidHS_ln1 ( ),
	. RxActiveHS_ln1 ( ),
	. RxSyncHS_ln1 ( ),
	. ext_TxDataHS_ln2 ( )
,
	. ext_TxRequestHS_ln2 ( ),
	. TxReadyHS_ln2 ( ),
	. ext_Enable_ln2 ( ),
	. ext_TxRequestEsc_ln2 ( ),
	. ext_TxUlpsEsc_ln2 ( ),
	. ext_TxLpdtEsc_ln2 ( ),
	. ext_TxUlpsExit_ln2 ( ),
	. TxReadyEsc_ln2 ( ),
	. ext_TxTriggerEsc_ln2 ( )
,
	. ext_TxDataEsc_ln2 ( )
,
	. ext_TxValidEsc_ln2 ( ),
	. ext_ForceTxStopmode_ln2 ( ),
	. ext_TurnRequest_ln2 ( ),
	. ext_TurnDisable_ln2 ( ),
	. ext_ForceRxmode_ln2 ( ),
	. RxClkEsc_ln2 ( ),
	. RxLpdtEsc_ln2 ( ),
	. RxUlpsEsc_ln2 ( ),
	. RxTriggerEsc_ln2 ( )
,
	. RxDataEsc_ln2 ( )
,
	. RxValidEsc_ln2 ( ),
	. Direction_ln2 ( ),
	. Stopstate_ln2 ( ),
	. UlpsActiveNot_ln2 ( ),
	. ErrSotHS_ln2 ( ),
	. ErrSotSyncHS_ln2 ( ),
	. ErrEsc_ln2 ( ),
	. ErrSyncEsc_ln2 ( ),
	. ErrControl_ln2 ( ),
	. ErrContentionLp0_ln2 ( ),
	. ErrContentionLp1_ln2 ( ),
	. RxDataHS_ln2 ( )
,
	. RxValidHS_ln2 ( ),
	. RxActiveHS_ln2 ( ),
	. RxSyncHS_ln2 ( ),
	. ext_TxDataHS_ln3 ( )
,
	. ext_TxRequestHS_ln3 ( ),
	. TxReadyHS_ln3 ( ),
	. ext_Enable_ln3 ( ),
	. ext_TxRequestEsc_ln3 ( ),
	. ext_TxUlpsEsc_ln3 ( ),
	. ext_TxLpdtEsc_ln3 ( ),
	. ext_TxUlpsExit_ln3 ( ),
	. TxReadyEsc_ln3 ( ),
	. ext_TxTriggerEsc_ln3 ( )
,
	. ext_TxDataEsc_ln3 ( )
,
	. ext_TxValidEsc_ln3 ( ),
	. ext_ForceTxStopmode_ln3 ( ),
	. ext_TurnRequest_ln3 ( ),
	. ext_TurnDisable_ln3 ( ),
	. ext_ForceRxmode_ln3 ( ),
	. RxClkEsc_ln3 ( ),
	. RxLpdtEsc_ln3 ( ),
	. RxUlpsEsc_ln3 ( ),
	. RxTriggerEsc_ln3 ( )
,
	. RxDataEsc_ln3 ( )
,
	. RxValidEsc_ln3 ( ),
	. Direction_ln3 ( ),
	. Stopstate_ln3 ( ),
	. UlpsActiveNot_ln3 ( ),
	. ErrSotHS_ln3 ( ),
	. ErrSotSyncHS_ln3 ( ),
	. ErrEsc_ln3 ( ),
	. ErrSyncEsc_ln3 ( ),
	. ErrControl_ln3 ( ),
	. ErrContentionLp0_ln3 ( ),
	. ErrContentionLp1_ln3 ( ),
	. RxDataHS_ln3 ( )
,
	. RxValidHS_ln3 ( ),
	. RxActiveHS_ln3 ( ),
	. RxSyncHS_ln3 ( ),
	. tx_dphy_rdy ( \mipi_inst_u_mipi1|tx_dphy_rdy_net  )
);
defparam mipi_inst_u_mipi1.HSEL = 0;
defparam mipi_inst_u_mipi1.PLACE_LOCATION = "C2R8.mipi_wrap.mipi1_top";
defparam mipi_inst_u_mipi1.RX_RCAL_OVRD = 0;
defparam mipi_inst_u_mipi1.RCAL_SEL = 0;
defparam mipi_inst_u_mipi1.PCK_LOCATION = "NONE";
defparam mipi_inst_u_mipi1.DELAY_BUF_NUM = 0;
defparam mipi_inst_u_mipi1.CLK_DLY = 0;
defparam mipi_inst_u_mipi1.DSI_CSI = 1;
defparam mipi_inst_u_mipi1.mipi_sel = "0";
defparam mipi_inst_u_mipi1.EXT_PPI_EN = 0;
defparam mipi_inst_u_mipi1.TX_RCAL_OVRD = 0;
LUT6 ii2615 (
	. xy ( \ii2615|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2615.PLACE_LOCATION = "C10R9.le_tile.le_guts.lp0.lut_0";
defparam ii2615.PCK_LOCATION = "C10R9.lp0.lut_0";
defparam ii2615.config_data = 64'b1111010111100100101100011010000011110101111001001011000110100000;
REG \mcu_arbiter_u_psram_dsel_reg[1]  (
	. qx ( \mcu_arbiter_u_psram_dsel_reg[1]|qx_net  ),
	. di ( \u_8051_u_h6_8051|memaddr_comb[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam \mcu_arbiter_u_psram_dsel_reg[1] .latch_mode = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .init = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .PLACE_LOCATION = "C16R26.le_tile.le_guts.lp0.reg0";
defparam \mcu_arbiter_u_psram_dsel_reg[1] .sr_inv = 1;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .sync_mode = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .no_sr = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .sr_value = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .PCK_LOCATION = "C16R26.lp0.reg0";
defparam \mcu_arbiter_u_psram_dsel_reg[1] .clk_inv = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .en_inv = 0;
defparam \mcu_arbiter_u_psram_dsel_reg[1] .always_en = 1;
MIPI_TOP mipi_inst_u_mipi2 (
	. CN ( {
		/* CN [4] */ \mipi_inst_u_mipi2|CN[4]_net ,
		/* CN [3] */ \mipi_inst_u_mipi2|CN[3]_net ,
		/* CN [2] */ \mipi_inst_u_mipi2|CN[2]_net ,
		/* CN [1] */ \mipi_inst_u_mipi2|CN[1]_net ,
		/* CN [0] */ \mipi_inst_u_mipi2|CN[0]_net 
	} ),
	. CM ( {
		/* CM [7] */ \mipi_inst_u_mipi2|CM[7]_net ,
		/* CM [6] */ \mipi_inst_u_mipi2|CM[6]_net ,
		/* CM [5] */ \mipi_inst_u_mipi2|CM[5]_net ,
		/* CM [4] */ \mipi_inst_u_mipi2|CM[4]_net ,
		/* CM [3] */ \mipi_inst_u_mipi2|CM[3]_net ,
		/* CM [2] */ \mipi_inst_u_mipi2|CM[2]_net ,
		/* CM [1] */ \mipi_inst_u_mipi2|CM[1]_net ,
		/* CM [0] */ \mipi_inst_u_mipi2|CM[0]_net 
	} ),
	. CO ( {
		/* CO [1] */ \mipi_inst_u_mipi2|CO[1]_net ,
		/* CO [0] */ \mipi_inst_u_mipi2|CO[0]_net 
	} ),
	. port_sel ( {
		/* port_sel [1] */ \GND_0_inst|Y_net ,
		/* port_sel [0] */ \VCC_0_inst|Y_net 
	} ),
	. enable_raw_dsi_port ( \VCC_0_inst|Y_net  ),
	. enable_dpi_port ( \GND_0_inst|Y_net  ),
	. TxEscClk ( \u_pll_pll_u0|CO1_net  ),
	. RxEscClk ( \u_pll_pll_u0|CO1_net  ),
	. reset_n ( \ii2048|xy_net  ),
	. reset_esc_n ( \ii2048|xy_net  ),
	. clk_periph ( ),
	. RxSyncHS ( ),
	. RxActiveHS ( ),
	. RxLpdtEsc ( ),
	. periph_dpi_vsync ( ),
	. periph_dpi_hsync ( ),
	. periph_dpi_de ( ),
	. periph_dpi_d ( )
,
	. periph_dpi_sd ( ),
	. periph_dpi_cm ( ),
	. periph_dpi_peripheral_output_dropped ( ),
	. periph_rx_cmd ( )
,
	. periph_rx_cmd_valid ( ),
	. periph_rx_payload ( )
,
	. periph_rx_payload_valid ( ),
	. periph_rx_payload_valid_last ( ),
	. periph_rx_trigger ( )
,
	. periph_rx_trigger_valid ( ),
	. periph_ecc_one_bit_err ( ),
	. periph_ecc_two_bit_err ( ),
	. periph_ecc_one_bit_err_pos ( )
,
	. periph_ecc_err ( ),
	. periph_ecc_err_pos ( )
,
	. periph_crc_err ( ),
	. periph_te_enable ( ),
	. periph_te_rdy ( ),
	. periph_te_ack ( ),
	. periph_te_event_in ( ),
	. periph_te_fail ( ),
	. periph_rx_ulps_active ( )
,
	. periph_rx_ulps_mark_active ( )
,
	. periph_tx_payload ( )
,
	. periph_tx_payload_en ( ),
	. periph_tx_payload_en_last ( ),
	. periph_tx_cmd_vc ( )
,
	. periph_tx_cmd_data_type ( )
,
	. periph_tx_cmd_byte_count ( )
,
	. periph_tx_cmd_req ( ),
	. periph_tx_cmd_ack ( ),
	. periph_tx_timeout_error ( ),
	. periph_trigger_req ( ),
	. periph_trigger_ack ( ),
	. periph_trigger_send ( )
,
	. periph_dphy_direction ( ),
	. hs_rx_timeout ( ),
	. lp_tx_timeout ( ),
	. periph_bta_timeout ( ),
	. dpi_pclk ( ),
	. reset_dpi_n ( ),
	. host_dpi_vsync ( ),
	. host_dpi_hsync ( ),
	. host_dpi_de ( ),
	. host_dpi_d ( )
,
	. host_dpi_sd ( ),
	. host_dpi_cm ( ),
	. dpi_host_underrun_err ( ),
	. host_tx_cmd_vc ( {
		/* host_tx_cmd_vc [1] */ \ii2078|xy_net ,
		/* host_tx_cmd_vc [0] */ \ii2077|xy_net 
	} ),
	. host_tx_cmd_data_type ( {
		/* host_tx_cmd_data_type [5] */ \ii2073|xy_net ,
		/* host_tx_cmd_data_type [4] */ \ii2072|xy_net ,
		/* host_tx_cmd_data_type [3] */ \ii2071|xy_net ,
		/* host_tx_cmd_data_type [2] */ \ii2070|xy_net ,
		/* host_tx_cmd_data_type [1] */ \ii2069|xy_net ,
		/* host_tx_cmd_data_type [0] */ \ii2068|xy_net 
	} ),
	. host_tx_cmd_byte_count ( {
		/* host_tx_cmd_byte_count [15] */ \ii2058|xy_net ,
		/* host_tx_cmd_byte_count [14] */ \ii2057|xy_net ,
		/* host_tx_cmd_byte_count [13] */ \ii2056|xy_net ,
		/* host_tx_cmd_byte_count [12] */ \ii2055|xy_net ,
		/* host_tx_cmd_byte_count [11] */ \ii2054|xy_net ,
		/* host_tx_cmd_byte_count [10] */ \ii2053|xy_net ,
		/* host_tx_cmd_byte_count [9] */ \ii2067|xy_net ,
		/* host_tx_cmd_byte_count [8] */ \ii2066|xy_net ,
		/* host_tx_cmd_byte_count [7] */ \ii2065|xy_net ,
		/* host_tx_cmd_byte_count [6] */ \ii2064|xy_net ,
		/* host_tx_cmd_byte_count [5] */ \ii2063|xy_net ,
		/* host_tx_cmd_byte_count [4] */ \ii2062|xy_net ,
		/* host_tx_cmd_byte_count [3] */ \ii2061|xy_net ,
		/* host_tx_cmd_byte_count [2] */ \ii2060|xy_net ,
		/* host_tx_cmd_byte_count [1] */ \ii2059|xy_net ,
		/* host_tx_cmd_byte_count [0] */ \ii2052|xy_net 
	} ),
	. host_tx_cmd_ack ( \mipi_inst_u_mipi2|host_tx_cmd_ack_net  ),
	. host_tx_cmd_req ( \ii2076|xy_net  ),
	. host_tx_payload ( {
		/* host_tx_payload [31] */ \ii2104|xy_net ,
		/* host_tx_payload [30] */ \ii2103|xy_net ,
		/* host_tx_payload [29] */ \ii2101|xy_net ,
		/* host_tx_payload [28] */ \ii2100|xy_net ,
		/* host_tx_payload [27] */ \ii2099|xy_net ,
		/* host_tx_payload [26] */ \ii2098|xy_net ,
		/* host_tx_payload [25] */ \ii2097|xy_net ,
		/* host_tx_payload [24] */ \ii2096|xy_net ,
		/* host_tx_payload [23] */ \ii2095|xy_net ,
		/* host_tx_payload [22] */ \ii2094|xy_net ,
		/* host_tx_payload [21] */ \ii2093|xy_net ,
		/* host_tx_payload [20] */ \ii2092|xy_net ,
		/* host_tx_payload [19] */ \ii2090|xy_net ,
		/* host_tx_payload [18] */ \ii2089|xy_net ,
		/* host_tx_payload [17] */ \ii2088|xy_net ,
		/* host_tx_payload [16] */ \ii2087|xy_net ,
		/* host_tx_payload [15] */ \ii2086|xy_net ,
		/* host_tx_payload [14] */ \ii2085|xy_net ,
		/* host_tx_payload [13] */ \ii2084|xy_net ,
		/* host_tx_payload [12] */ \ii2083|xy_net ,
		/* host_tx_payload [11] */ \ii2082|xy_net ,
		/* host_tx_payload [10] */ \ii2081|xy_net ,
		/* host_tx_payload [9] */ \ii2111|xy_net ,
		/* host_tx_payload [8] */ \ii2110|xy_net ,
		/* host_tx_payload [7] */ \ii2109|xy_net ,
		/* host_tx_payload [6] */ \ii2108|xy_net ,
		/* host_tx_payload [5] */ \ii2107|xy_net ,
		/* host_tx_payload [4] */ \ii2106|xy_net ,
		/* host_tx_payload [3] */ \ii2105|xy_net ,
		/* host_tx_payload [2] */ \ii2102|xy_net ,
		/* host_tx_payload [1] */ \ii2091|xy_net ,
		/* host_tx_payload [0] */ \ii2080|xy_net 
	} ),
	. host_tx_payload_en ( \mipi_inst_u_mipi2|host_tx_payload_en_net  ),
	. host_tx_payload_en_last ( \mipi_inst_u_mipi2|host_tx_payload_en_last_net  ),
	. host_tx_hs_mode ( \ii2079|xy_net  ),
	. host_tx_active ( \mipi_inst_u_mipi2|host_tx_active_net  ),
	. host_tx_ulps_enable ( {
		/* host_tx_ulps_enable [4] */ \GND_0_inst|Y_net ,
		/* host_tx_ulps_enable [3] */ \GND_0_inst|Y_net ,
		/* host_tx_ulps_enable [2] */ \GND_0_inst|Y_net ,
		/* host_tx_ulps_enable [1] */ \GND_0_inst|Y_net ,
		/* host_tx_ulps_enable [0] */ \GND_0_inst|Y_net 
	} ),
	. host_tx_ulps_active ( )
,
	. host_dphy_turnaround ( \GND_0_inst|Y_net  ),
	. host_dphy_direction ( ),
	. host_trigger_req ( \GND_0_inst|Y_net  ),
	. host_trigger_send ( {
		/* host_trigger_send [1] */ \GND_0_inst|Y_net ,
		/* host_trigger_send [0] */ \GND_0_inst|Y_net 
	} ),
	. host_trigger_ack ( ),
	. host_rx_payload ( )
,
	. host_rx_payload_valid ( ),
	. host_rx_payload_valid_last ( ),
	. host_rx_cmd_valid ( ),
	. host_rx_cmd_vc ( )
,
	. host_rx_cmd_data_type ( )
,
	. host_rx_cmd_byte_count ( )
,
	. host_ecc_one_bit_err ( ),
	. host_ecc_two_bit_err ( ),
	. host_ecc_one_bit_err_pos ( )
,
	. host_ecc_err ( ),
	. host_ecc_err_pos ( )
,
	. host_crc_err ( ),
	. host_hs_tx_timeout ( ),
	. host_lp_rx_timeout ( ),
	. host_bta_timeout ( ),
	. pclk_reset_n ( \ii1982|xy_net  ),
	. pclk ( \u_pll_pll_u0|CO3_net  ),
	. paddr ( {
		/* paddr [17] */ \GND_0_inst|Y_net ,
		/* paddr [16] */ \GND_0_inst|Y_net ,
		/* paddr [15] */ \GND_0_inst|Y_net ,
		/* paddr [14] */ \GND_0_inst|Y_net ,
		/* paddr [13] */ \GND_0_inst|Y_net ,
		/* paddr [12] */ \GND_0_inst|Y_net ,
		/* paddr [11] */ \GND_0_inst|Y_net ,
		/* paddr [10] */ \GND_0_inst|Y_net ,
		/* paddr [9] */ \u_8051_u_h6_8051|memaddr_comb[9]_net ,
		/* paddr [8] */ \u_8051_u_h6_8051|memaddr_comb[8]_net ,
		/* paddr [7] */ \u_8051_u_h6_8051|memaddr_comb[7]_net ,
		/* paddr [6] */ \u_8051_u_h6_8051|memaddr_comb[6]_net ,
		/* paddr [5] */ \u_8051_u_h6_8051|memaddr_comb[5]_net ,
		/* paddr [4] */ \u_8051_u_h6_8051|memaddr_comb[4]_net ,
		/* paddr [3] */ \u_8051_u_h6_8051|memaddr_comb[3]_net ,
		/* paddr [2] */ \u_8051_u_h6_8051|memaddr_comb[2]_net ,
		/* paddr [1] */ \GND_0_inst|Y_net ,
		/* paddr [0] */ \GND_0_inst|Y_net 
	} ),
	. pwrite ( \mcu_arbiter_u_emif2apb_u0_dbuf_u_delaybuf|xy_net  ),
	. psel ( \ii2112|xy_net  ),
	. penable ( \ii2050|xy_net  ),
	. pwdata ( {
		/* pwdata [31] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_31__u_delaybuf|xy_net ,
		/* pwdata [30] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_30__u_delaybuf|xy_net ,
		/* pwdata [29] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_29__u_delaybuf|xy_net ,
		/* pwdata [28] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_28__u_delaybuf|xy_net ,
		/* pwdata [27] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_27__u_delaybuf|xy_net ,
		/* pwdata [26] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_26__u_delaybuf|xy_net ,
		/* pwdata [25] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_25__u_delaybuf|xy_net ,
		/* pwdata [24] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_24__u_delaybuf|xy_net ,
		/* pwdata [23] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_23__u_delaybuf|xy_net ,
		/* pwdata [22] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_22__u_delaybuf|xy_net ,
		/* pwdata [21] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_21__u_delaybuf|xy_net ,
		/* pwdata [20] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_20__u_delaybuf|xy_net ,
		/* pwdata [19] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_19__u_delaybuf|xy_net ,
		/* pwdata [18] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_18__u_delaybuf|xy_net ,
		/* pwdata [17] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_17__u_delaybuf|xy_net ,
		/* pwdata [16] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_16__u_delaybuf|xy_net ,
		/* pwdata [15] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_15__u_delaybuf|xy_net ,
		/* pwdata [14] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_14__u_delaybuf|xy_net ,
		/* pwdata [13] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_13__u_delaybuf|xy_net ,
		/* pwdata [12] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_12__u_delaybuf|xy_net ,
		/* pwdata [11] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_11__u_delaybuf|xy_net ,
		/* pwdata [10] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_10__u_delaybuf|xy_net ,
		/* pwdata [9] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_9__u_delaybuf|xy_net ,
		/* pwdata [8] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_8__u_delaybuf|xy_net ,
		/* pwdata [7] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_7__u_delaybuf|xy_net ,
		/* pwdata [6] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_6__u_delaybuf|xy_net ,
		/* pwdata [5] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_5__u_delaybuf|xy_net ,
		/* pwdata [4] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_4__u_delaybuf|xy_net ,
		/* pwdata [3] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_3__u_delaybuf|xy_net ,
		/* pwdata [2] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_2__u_delaybuf|xy_net ,
		/* pwdata [1] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_1__u_delaybuf|xy_net ,
		/* pwdata [0] */ \mcu_arbiter_u_emif2apb_u0_dx32_genblk1_0__u_delaybuf|xy_net 
	} ),
	. prdata ( {
		/* prdata [31] */ \mipi_inst_u_mipi2|prdata[31]_net ,
		/* prdata [30] */ \mipi_inst_u_mipi2|prdata[30]_net ,
		/* prdata [29] */ \mipi_inst_u_mipi2|prdata[29]_net ,
		/* prdata [28] */ \mipi_inst_u_mipi2|prdata[28]_net ,
		/* prdata [27] */ \mipi_inst_u_mipi2|prdata[27]_net ,
		/* prdata [26] */ \mipi_inst_u_mipi2|prdata[26]_net ,
		/* prdata [25] */ \mipi_inst_u_mipi2|prdata[25]_net ,
		/* prdata [24] */ \mipi_inst_u_mipi2|prdata[24]_net ,
		/* prdata [23] */ \mipi_inst_u_mipi2|prdata[23]_net ,
		/* prdata [22] */ \mipi_inst_u_mipi2|prdata[22]_net ,
		/* prdata [21] */ \mipi_inst_u_mipi2|prdata[21]_net ,
		/* prdata [20] */ \mipi_inst_u_mipi2|prdata[20]_net ,
		/* prdata [19] */ \mipi_inst_u_mipi2|prdata[19]_net ,
		/* prdata [18] */ \mipi_inst_u_mipi2|prdata[18]_net ,
		/* prdata [17] */ \mipi_inst_u_mipi2|prdata[17]_net ,
		/* prdata [16] */ \mipi_inst_u_mipi2|prdata[16]_net ,
		/* prdata [15] */ \mipi_inst_u_mipi2|prdata[15]_net ,
		/* prdata [14] */ \mipi_inst_u_mipi2|prdata[14]_net ,
		/* prdata [13] */ \mipi_inst_u_mipi2|prdata[13]_net ,
		/* prdata [12] */ \mipi_inst_u_mipi2|prdata[12]_net ,
		/* prdata [11] */ \mipi_inst_u_mipi2|prdata[11]_net ,
		/* prdata [10] */ \mipi_inst_u_mipi2|prdata[10]_net ,
		/* prdata [9] */ \mipi_inst_u_mipi2|prdata[9]_net ,
		/* prdata [8] */ \mipi_inst_u_mipi2|prdata[8]_net ,
		/* prdata [7] */ \mipi_inst_u_mipi2|prdata[7]_net ,
		/* prdata [6] */ \mipi_inst_u_mipi2|prdata[6]_net ,
		/* prdata [5] */ \mipi_inst_u_mipi2|prdata[5]_net ,
		/* prdata [4] */ \mipi_inst_u_mipi2|prdata[4]_net ,
		/* prdata [3] */ \mipi_inst_u_mipi2|prdata[3]_net ,
		/* prdata [2] */ \mipi_inst_u_mipi2|prdata[2]_net ,
		/* prdata [1] */ \mipi_inst_u_mipi2|prdata[1]_net ,
		/* prdata [0] */ \mipi_inst_u_mipi2|prdata[0]_net 
	} ),
	. pready ( \mipi_inst_u_mipi2|pready_net  ),
	. clk ( \mipi_inst_u_mipi2|clk_net  ),
	. RxByteClkHS ( ),
	. CLKP ( ),
	. CLKN ( ),
	. DATAN0 ( ),
	. DATAP0 ( ),
	. DATAN1 ( ),
	. DATAP1 ( ),
	. DATAN2 ( ),
	. DATAP2 ( ),
	. DATAN3 ( ),
	. DATAP3 ( ),
	. LOCK ( \mipi_inst_u_mipi_pll|LOCK_net  ),
	. BITCLK ( \mipi_inst_u_mipi_pll|CLKOUT2_net  ),
	. PD_DPHY ( \ii2049|xy_net  ),
	. ENP_DESER ( \GND_0_inst|Y_net  ),
	. TEST_ENBL ( {
		/* TEST_ENBL [5] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [4] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [3] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [2] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [1] */ \GND_0_inst|Y_net ,
		/* TEST_ENBL [0] */ \GND_0_inst|Y_net 
	} ),
	. TEST_PATTERN ( )
,
	. D0_LB_PASS ( )
,
	. D1_LB_PASS ( )
,
	. D2_LB_PASS ( )
,
	. D3_LB_PASS ( )
,
	. D0_LB_ERR_CNT ( )
,
	. D1_LB_ERR_CNT ( )
,
	. D2_LB_ERR_CNT ( )
,
	. D3_LB_ERR_CNT ( )
,
	. D0_LB_BYTE_CNT ( )
,
	. D1_LB_BYTE_CNT ( )
,
	. D2_LB_BYTE_CNT ( )
,
	. D3_LB_BYTE_CNT ( )
,
	. D0_LB_ACTIVE ( )
,
	. D1_LB_ACTIVE ( )
,
	. D2_LB_ACTIVE ( )
,
	. D3_LB_ACTIVE ( )
,
	. D0_LB_VALID ( )
,
	. D1_LB_VALID ( )
,
	. D2_LB_VALID ( )
,
	. D3_LB_VALID ( )
,
	. CLK_LB_ACTIVE ( ),
	. DC_TEST_OUT ( )
,
	. AUTO_PD_EN ( \GND_0_inst|Y_net  ),
	. ext_TxRequestHS_lnclk ( ),
	. Stopstate_lnclk ( ),
	. ext_TxUlpsClk_lnclk ( ),
	. ext_TxUlpsExit_lnclk ( ),
	. UlpsActiveNot_lnclk ( ),
	. RxUlpsClkNot ( ),
	. RxClkActiveHS ( ),
	. ext_Enable_lnclk ( ),
	. ext_TxDataHS_ln0 ( )
,
	. ext_TxRequestHS_ln0 ( ),
	. TxReadyHS_ln0 ( ),
	. ext_Enable_ln0 ( ),
	. ext_TxRequestEsc_ln0 ( ),
	. ext_TxUlpsEsc_ln0 ( ),
	. ext_TxLpdtEsc_ln0 ( ),
	. ext_TxUlpsExit_ln0 ( ),
	. TxReadyEsc_ln0 ( ),
	. ext_TxTriggerEsc_ln0 ( )
,
	. ext_TxDataEsc_ln0 ( )
,
	. ext_TxValidEsc_ln0 ( ),
	. ext_ForceTxStopmode_ln0 ( ),
	. ext_TurnRequest_ln0 ( ),
	. ext_TurnDisable_ln0 ( ),
	. ext_ForceRxmode_ln0 ( ),
	. RxClkEsc_ln0 ( ),
	. RxLpdtEsc_ln0 ( ),
	. RxUlpsEsc_ln0 ( ),
	. RxTriggerEsc_ln0 ( )
,
	. RxDataEsc_ln0 ( )
,
	. RxValidEsc_ln0 ( ),
	. Direction_ln0 ( ),
	. Stopstate_ln0 ( ),
	. UlpsActiveNot_ln0 ( ),
	. ErrSotHS_ln0 ( ),
	. ErrSotSyncHS_ln0 ( ),
	. ErrEsc_ln0 ( ),
	. ErrSyncEsc_ln0 ( ),
	. ErrControl_ln0 ( ),
	. ErrContentionLp0_ln0 ( ),
	. ErrContentionLp1_ln0 ( ),
	. RxDataHS_ln0 ( )
,
	. RxValidHS_ln0 ( ),
	. RxActiveHS_ln0 ( ),
	. RxSyncHS_ln0 ( ),
	. ext_TxDataHS_ln1 ( )
,
	. ext_TxRequestHS_ln1 ( ),
	. TxReadyHS_ln1 ( ),
	. ext_Enable_ln1 ( ),
	. ext_TxRequestEsc_ln1 ( ),
	. ext_TxUlpsEsc_ln1 ( ),
	. ext_TxLpdtEsc_ln1 ( ),
	. ext_TxUlpsExit_ln1 ( ),
	. TxReadyEsc_ln1 ( ),
	. ext_TxTriggerEsc_ln1 ( )
,
	. ext_TxDataEsc_ln1 ( )
,
	. ext_TxValidEsc_ln1 ( ),
	. ext_ForceTxStopmode_ln1 ( ),
	. ext_TurnRequest_ln1 ( ),
	. ext_TurnDisable_ln1 ( ),
	. ext_ForceRxmode_ln1 ( ),
	. RxClkEsc_ln1 ( ),
	. RxLpdtEsc_ln1 ( ),
	. RxUlpsEsc_ln1 ( ),
	. RxTriggerEsc_ln1 ( )
,
	. RxDataEsc_ln1 ( )
,
	. RxValidEsc_ln1 ( ),
	. Direction_ln1 ( ),
	. Stopstate_ln1 ( ),
	. UlpsActiveNot_ln1 ( ),
	. ErrSotHS_ln1 ( ),
	. ErrSotSyncHS_ln1 ( ),
	. ErrEsc_ln1 ( ),
	. ErrSyncEsc_ln1 ( ),
	. ErrControl_ln1 ( ),
	. ErrContentionLp0_ln1 ( ),
	. ErrContentionLp1_ln1 ( ),
	. RxDataHS_ln1 ( )
,
	. RxValidHS_ln1 ( ),
	. RxActiveHS_ln1 ( ),
	. RxSyncHS_ln1 ( ),
	. ext_TxDataHS_ln2 ( )
,
	. ext_TxRequestHS_ln2 ( ),
	. TxReadyHS_ln2 ( ),
	. ext_Enable_ln2 ( ),
	. ext_TxRequestEsc_ln2 ( ),
	. ext_TxUlpsEsc_ln2 ( ),
	. ext_TxLpdtEsc_ln2 ( ),
	. ext_TxUlpsExit_ln2 ( ),
	. TxReadyEsc_ln2 ( ),
	. ext_TxTriggerEsc_ln2 ( )
,
	. ext_TxDataEsc_ln2 ( )
,
	. ext_TxValidEsc_ln2 ( ),
	. ext_ForceTxStopmode_ln2 ( ),
	. ext_TurnRequest_ln2 ( ),
	. ext_TurnDisable_ln2 ( ),
	. ext_ForceRxmode_ln2 ( ),
	. RxClkEsc_ln2 ( ),
	. RxLpdtEsc_ln2 ( ),
	. RxUlpsEsc_ln2 ( ),
	. RxTriggerEsc_ln2 ( )
,
	. RxDataEsc_ln2 ( )
,
	. RxValidEsc_ln2 ( ),
	. Direction_ln2 ( ),
	. Stopstate_ln2 ( ),
	. UlpsActiveNot_ln2 ( ),
	. ErrSotHS_ln2 ( ),
	. ErrSotSyncHS_ln2 ( ),
	. ErrEsc_ln2 ( ),
	. ErrSyncEsc_ln2 ( ),
	. ErrControl_ln2 ( ),
	. ErrContentionLp0_ln2 ( ),
	. ErrContentionLp1_ln2 ( ),
	. RxDataHS_ln2 ( )
,
	. RxValidHS_ln2 ( ),
	. RxActiveHS_ln2 ( ),
	. RxSyncHS_ln2 ( ),
	. ext_TxDataHS_ln3 ( )
,
	. ext_TxRequestHS_ln3 ( ),
	. TxReadyHS_ln3 ( ),
	. ext_Enable_ln3 ( ),
	. ext_TxRequestEsc_ln3 ( ),
	. ext_TxUlpsEsc_ln3 ( ),
	. ext_TxLpdtEsc_ln3 ( ),
	. ext_TxUlpsExit_ln3 ( ),
	. TxReadyEsc_ln3 ( ),
	. ext_TxTriggerEsc_ln3 ( )
,
	. ext_TxDataEsc_ln3 ( )
,
	. ext_TxValidEsc_ln3 ( ),
	. ext_ForceTxStopmode_ln3 ( ),
	. ext_TurnRequest_ln3 ( ),
	. ext_TurnDisable_ln3 ( ),
	. ext_ForceRxmode_ln3 ( ),
	. RxClkEsc_ln3 ( ),
	. RxLpdtEsc_ln3 ( ),
	. RxUlpsEsc_ln3 ( ),
	. RxTriggerEsc_ln3 ( )
,
	. RxDataEsc_ln3 ( )
,
	. RxValidEsc_ln3 ( ),
	. Direction_ln3 ( ),
	. Stopstate_ln3 ( ),
	. UlpsActiveNot_ln3 ( ),
	. ErrSotHS_ln3 ( ),
	. ErrSotSyncHS_ln3 ( ),
	. ErrEsc_ln3 ( ),
	. ErrSyncEsc_ln3 ( ),
	. ErrControl_ln3 ( ),
	. ErrContentionLp0_ln3 ( ),
	. ErrContentionLp1_ln3 ( ),
	. RxDataHS_ln3 ( )
,
	. RxValidHS_ln3 ( ),
	. RxActiveHS_ln3 ( ),
	. RxSyncHS_ln3 ( ),
	. tx_dphy_rdy ( \mipi_inst_u_mipi2|tx_dphy_rdy_net  )
);
defparam mipi_inst_u_mipi2.HSEL = 0;
defparam mipi_inst_u_mipi2.PLACE_LOCATION = "C2R24.mipi_wrap.mipi2_top";
defparam mipi_inst_u_mipi2.RX_RCAL_OVRD = 0;
defparam mipi_inst_u_mipi2.RCAL_SEL = 0;
defparam mipi_inst_u_mipi2.PCK_LOCATION = "NONE";
defparam mipi_inst_u_mipi2.DELAY_BUF_NUM = 0;
defparam mipi_inst_u_mipi2.CLK_DLY = 1;
defparam mipi_inst_u_mipi2.DSI_CSI = 1;
defparam mipi_inst_u_mipi2.mipi_sel = "1";
defparam mipi_inst_u_mipi2.EXT_PPI_EN = 0;
defparam mipi_inst_u_mipi2.TX_RCAL_OVRD = 0;
LUT6 ii2616 (
	. xy ( \ii2616|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[2]|qx_net  )
);
defparam ii2616.PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.lut_0";
defparam ii2616.PCK_LOCATION = "C14R9.lp0.lut_0";
defparam ii2616.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12]|qx_net  ),
	. di ( \ii2871|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[12] .always_en = 1;
LUT6 ii2617 (
	. xy ( \ii2617|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2616|xy_net  ),
	. f1 ( \ii2615|xy_net  ),
	. f0 ( \ii2614|xy_net  )
);
defparam ii2617.PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.lut_0";
defparam ii2617.PCK_LOCATION = "C14R8.lp0.lut_0";
defparam ii2617.config_data = 64'b1111000010101010110011001100110011110000101010101100110011001100;
REG glue_rd_cmd_flag_reg (
	. qx ( \glue_rd_cmd_flag_reg|qx_net  ),
	. di ( \ii2137|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rd_cmd_flag_reg.latch_mode = 0;
defparam glue_rd_cmd_flag_reg.init = 0;
defparam glue_rd_cmd_flag_reg.PLACE_LOCATION = "C14R24.le_tile.le_guts.lp0.reg0";
defparam glue_rd_cmd_flag_reg.sr_inv = 1;
defparam glue_rd_cmd_flag_reg.sync_mode = 0;
defparam glue_rd_cmd_flag_reg.no_sr = 0;
defparam glue_rd_cmd_flag_reg.sr_value = 0;
defparam glue_rd_cmd_flag_reg.PCK_LOCATION = "C14R24.lp0.reg0";
defparam glue_rd_cmd_flag_reg.clk_inv = 0;
defparam glue_rd_cmd_flag_reg.en_inv = 0;
defparam glue_rd_cmd_flag_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4]|qx_net  ),
	. di ( \ii2917|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[4] .always_en = 1;
LUT6 ii2618 (
	. xy ( \ii2618|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2618.PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.lut_0";
defparam ii2618.PCK_LOCATION = "C14R9.lp0.lut_0";
defparam ii2618.config_data = 64'b1111010111100100101100011010000011110101111001001011000110100000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[18] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[1] .always_en = 1;
LUT6 ii2619 (
	. xy ( \ii2619|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2619.PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.lut_0";
defparam ii2619.PCK_LOCATION = "C14R8.lp0.lut_0";
defparam ii2619.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2620 (
	. xy ( \ii2620|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[3]|qx_net  )
);
defparam ii2620.PLACE_LOCATION = "C14R9.le_tile.le_guts.lp0.lut_0";
defparam ii2620.PCK_LOCATION = "C14R9.lp0.lut_0";
defparam ii2620.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6]|qx_net  ),
	. di ( \ii2335|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[6] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. di ( \ii2656|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. di ( \ii2664|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20] .always_en = 1;
LUT6 ii2621 (
	. xy ( \ii2621|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2620|xy_net  ),
	. f1 ( \ii2619|xy_net  ),
	. f0 ( \ii2618|xy_net  )
);
defparam ii2621.PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.lut_0";
defparam ii2621.PCK_LOCATION = "C14R8.lp0.lut_0";
defparam ii2621.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5]|qx_net  ),
	. di ( \carry_9_7__ADD_5|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[5] .always_en = 1;
LUT6 ii2622 (
	. xy ( \ii2622|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2622.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2622.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2622.config_data = 64'b1111010111100100101100011010000011110101111001001011000110100000;
LUT6 ii2623 (
	. xy ( \ii2623|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2623.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2623.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2623.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2624 (
	. xy ( \ii2624|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[4]|qx_net  )
);
defparam ii2624.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2624.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2624.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
LUT6 ii2625 (
	. xy ( \ii2625|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2624|xy_net  ),
	. f1 ( \ii2623|xy_net  ),
	. f0 ( \ii2622|xy_net  )
);
defparam ii2625.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2625.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2625.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
LUT6 ii2626 (
	. xy ( \ii2626|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2626.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2626.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2626.config_data = 64'b1111010111100100101100011010000011110101111001001011000110100000;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13]|qx_net  ),
	. di ( \ii2873|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[13] .always_en = 1;
LUT6 ii2627 (
	. xy ( \ii2627|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2627.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2627.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2627.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5]|qx_net  ),
	. di ( \ii2919|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[5] .always_en = 1;
LUT6 ii2628 (
	. xy ( \ii2628|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[5]|qx_net  )
);
defparam ii2628.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2628.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2628.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[4]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[20] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[3]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .PLACE_LOCATION = "C14R27.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .PCK_LOCATION = "C14R27.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[19] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[2] .always_en = 1;
LUT6 ii2629 (
	. xy ( \ii2629|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2628|xy_net  ),
	. f1 ( \ii2627|xy_net  ),
	. f0 ( \ii2626|xy_net  )
);
defparam ii2629.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2629.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2629.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
LUT6 ii2630 (
	. xy ( \ii2630|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2630.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2630.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2630.config_data = 64'b1111010111100100101100011010000011110101111001001011000110100000;
REG glue_rx_packet_tx_packet_u_data_process_frame_start_reg (
	. qx ( \glue_rx_packet_tx_packet_u_data_process_frame_start_reg|qx_net  ),
	. di ( \ii2429|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.PCK_LOCATION = "C16R10.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_data_process_frame_start_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7]|qx_net  ),
	. di ( \ii2336|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .PLACE_LOCATION = "C8R4.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .PCK_LOCATION = "C8R4.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[7] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. di ( \ii2669|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21] .always_en = 1;
LUT6 ii2631 (
	. xy ( \ii2631|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2631.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2631.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2631.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG glue_pasm_tx_act_d_reg (
	. qx ( \glue_pasm_tx_act_d_reg|qx_net  ),
	. di ( \ii2136|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_pasm_tx_act_d_reg.latch_mode = 0;
defparam glue_pasm_tx_act_d_reg.init = 0;
defparam glue_pasm_tx_act_d_reg.PLACE_LOCATION = "C14R29.le_tile.le_guts.lp0.reg0";
defparam glue_pasm_tx_act_d_reg.sr_inv = 1;
defparam glue_pasm_tx_act_d_reg.sync_mode = 0;
defparam glue_pasm_tx_act_d_reg.no_sr = 0;
defparam glue_pasm_tx_act_d_reg.sr_value = 0;
defparam glue_pasm_tx_act_d_reg.PCK_LOCATION = "C14R29.lp0.reg0";
defparam glue_pasm_tx_act_d_reg.clk_inv = 0;
defparam glue_pasm_tx_act_d_reg.en_inv = 0;
defparam glue_pasm_tx_act_d_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6]|qx_net  ),
	. di ( \carry_9_7__ADD_6|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[6] .always_en = 1;
LUT6 ii2632 (
	. xy ( \ii2632|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[6]|qx_net  )
);
defparam ii2632.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2632.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2632.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
LUT6 ii2633 (
	. xy ( \ii2633|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2632|xy_net  ),
	. f1 ( \ii2631|xy_net  ),
	. f0 ( \ii2630|xy_net  )
);
defparam ii2633.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2633.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2633.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
LUT6 ii2634 (
	. xy ( \ii2634|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7]|qx_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2634.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2634.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2634.config_data = 64'b1111010111100100101100011010000011110101111001001011000110100000;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.PLACE_LOCATION = "C14R19.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.PCK_LOCATION = "C14R19.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_line_data_en_d_reg.always_en = 1;
LUT6 ii2635 (
	. xy ( \ii2635|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2635.PLACE_LOCATION = "C18R7.le_tile.le_guts.lp0.lut_0";
defparam ii2635.PCK_LOCATION = "C18R7.lp0.lut_0";
defparam ii2635.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
ADD1_A carry_9_5__ADD_0 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[0]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[0]|qx_net  ),
	. ci ( \VCC_0_inst|Y_net  ),
	. co ( \carry_9_5__ADD_0|co_net  ),
	. s ( \carry_9_5__ADD_0|s_net  )
);
defparam carry_9_5__ADD_0.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_0.a_inv = "true";
defparam carry_9_5__ADD_0.PCK_LOCATION = "C14R7.lp0.add2.add0";
LUT6 ii2636 (
	. xy ( \ii2636|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[7]|qx_net  )
);
defparam ii2636.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2636.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2636.config_data = 64'b1010101011110000111111111100110010101010111100000000000011001100;
ADD1_A carry_9_5__ADD_1 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[1]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[1]|qx_net  ),
	. ci ( \carry_9_5__ADD_0|co_net  ),
	. co ( \carry_9_5__ADD_1|co_net  ),
	. s ( \carry_9_5__ADD_1|s_net  )
);
defparam carry_9_5__ADD_1.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_1.a_inv = "true";
defparam carry_9_5__ADD_1.PCK_LOCATION = "C14R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14]|qx_net  ),
	. di ( \ii2875|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .PLACE_LOCATION = "C6R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .PCK_LOCATION = "C6R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[14] .always_en = 1;
LUT6 ii2637 (
	. xy ( \ii2637|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2636|xy_net  ),
	. f1 ( \ii2635|xy_net  ),
	. f0 ( \ii2634|xy_net  )
);
defparam ii2637.PLACE_LOCATION = "C18R8.le_tile.le_guts.lp0.lut_0";
defparam ii2637.PCK_LOCATION = "C18R8.lp0.lut_0";
defparam ii2637.config_data = 64'b1111000011001100101010101010101011110000110011001010101010101010;
ADD1_A carry_9_5__ADD_2 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[2]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[2]|qx_net  ),
	. ci ( \carry_9_5__ADD_1|co_net  ),
	. co ( \carry_9_5__ADD_2|co_net  ),
	. s ( \carry_9_5__ADD_2|s_net  )
);
defparam carry_9_5__ADD_2.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_2.a_inv = "true";
defparam carry_9_5__ADD_2.PCK_LOCATION = "C14R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6]|qx_net  ),
	. di ( \ii2921|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[6] .always_en = 1;
LUT6 ii2638 (
	. xy ( \ii2638|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f0 ( \ii2612|xy_net  )
);
defparam ii2638.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2638.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2638.config_data = 64'b0001000100110001000100110011001100010001001100010001001100110011;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[5]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[21] .always_en = 1;
ADD1_A carry_9_5__ADD_3 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[3]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[3]|qx_net  ),
	. ci ( \carry_9_5__ADD_2|co_net  ),
	. co ( \carry_9_5__ADD_3|co_net  ),
	. s ( \carry_9_5__ADD_3|s_net  )
);
defparam carry_9_5__ADD_3.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_3.a_inv = "true";
defparam carry_9_5__ADD_3.PCK_LOCATION = "C14R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[2] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[3]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[3] .always_en = 1;
LUT6 ii2639 (
	. xy ( \ii2639|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]|qx_net  )
);
defparam ii2639.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.lut_0";
defparam ii2639.PCK_LOCATION = "C18R11.lp0.lut_0";
defparam ii2639.config_data = 64'b0011010100000000001101010000111100110101111100000011010111111111;
LUT6 ii2640 (
	. xy ( \ii2640|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f1 ( \ii2639|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2640.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.lut_0";
defparam ii2640.PCK_LOCATION = "C18R12.lp0.lut_0";
defparam ii2640.config_data = 64'b1100000000000000110001010000000011001010000000001100111100000000;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8]|qx_net  ),
	. di ( \ii2337|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .PCK_LOCATION = "C10R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[8] .always_en = 0;
ADD1_A carry_9_5__ADD_4 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[4]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[4]|qx_net  ),
	. ci ( \carry_9_5__ADD_3|co_net  ),
	. co ( \carry_9_5__ADD_4|co_net  ),
	. s ( \carry_9_5__ADD_4|s_net  )
);
defparam carry_9_5__ADD_4.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_4.a_inv = "true";
defparam carry_9_5__ADD_4.PCK_LOCATION = "C14R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. di ( \ii2674|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22] .always_en = 1;
LUT6 ii2641 (
	. xy ( \ii2641|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[0]|qx_net  ),
	. f3 ( \ii2612|xy_net  ),
	. f2 ( \ii2582|xy_net  ),
	. f1 ( \ii2640|xy_net  ),
	. f0 ( \ii2638|xy_net  )
);
defparam ii2641.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.lut_0";
defparam ii2641.PCK_LOCATION = "C18R12.lp0.lut_0";
defparam ii2641.config_data = 64'b0001000100110011000100010001001100010001001100010001000100010001;
ADD1_A carry_9_5__ADD_5 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[5]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[5]|qx_net  ),
	. ci ( \carry_9_5__ADD_4|co_net  ),
	. co ( \carry_9_5__ADD_5|co_net  ),
	. s ( \carry_9_5__ADD_5|s_net  )
);
defparam carry_9_5__ADD_5.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_5.a_inv = "true";
defparam carry_9_5__ADD_5.PCK_LOCATION = "C14R7.lp0.add2.add0";
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7]|qx_net  ),
	. di ( \carry_9_7__ADD_7|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .PLACE_LOCATION = "C20R18.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .PCK_LOCATION = "C20R18.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[7] .always_en = 1;
REG glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg (
	. qx ( \glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg|qx_net  ),
	. di ( \ii3284|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.init = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.PLACE_LOCATION = "C14R17.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.PCK_LOCATION = "C14R17.lp0.reg0";
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_u_sync_delay_first_vs_delay_flag_reg.always_en = 1;
LUT6 ii2642 (
	. xy ( \ii2642|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]|qx_net  )
);
defparam ii2642.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.lut_0";
defparam ii2642.PCK_LOCATION = "C18R11.lp0.lut_0";
defparam ii2642.config_data = 64'b1100101011111111110010101111000011001010111111111100101011110000;
ADD1_A carry_9_5__ADD_6 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[6]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[6]|qx_net  ),
	. ci ( \carry_9_5__ADD_5|co_net  ),
	. co ( \carry_9_5__ADD_6|co_net  ),
	. s ( \carry_9_5__ADD_6|s_net  )
);
defparam carry_9_5__ADD_6.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_6.a_inv = "true";
defparam carry_9_5__ADD_6.PCK_LOCATION = "C14R7.lp0.add2.add0";
LUT6 ii2643 (
	. xy ( \ii2643|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \ii2642|xy_net  )
);
defparam ii2643.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2643.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2643.config_data = 64'b0101010100000000010111011111110001010101000000110101110111111111;
ADD1_A carry_9_5__ADD_7 (
	. a ( \glue_rx_packet_tx_packet_u_scaler_t8_out1_4_reg[7]|qx_net  ),
	. b ( \glue_rx_packet_tx_packet_u_scaler_t23_out1_reg[7]|qx_net  ),
	. ci ( \carry_9_5__ADD_6|co_net  ),
	. co ( \carry_9_5__ADD_7|co_net  ),
	. s ( \carry_9_5__ADD_7|s_net  )
);
defparam carry_9_5__ADD_7.PLACE_LOCATION = "C14R7.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_7.a_inv = "true";
defparam carry_9_5__ADD_7.PCK_LOCATION = "C14R7.lp0.add2.add0";
LUT6 ii2644 (
	. xy ( \ii2644|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[17]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]|qx_net  )
);
defparam ii2644.PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.lut_0";
defparam ii2644.PCK_LOCATION = "C16R12.lp0.lut_0";
defparam ii2644.config_data = 64'b0100000000000000011111110011001101000000000000000111111100110011;
ADD1_A carry_9_5__ADD_8 (
	. a ( \GND_0_inst|Y_net  ),
	. b ( \VCC_0_inst|Y_net  ),
	. ci ( \carry_9_5__ADD_7|co_net  ),
	. co ( \carry_9_5__ADD_8|co_net  ),
	. s ( )
);
defparam carry_9_5__ADD_8.PLACE_LOCATION = "C14R8.le_tile.le_guts.lp0.add2.add0";
defparam carry_9_5__ADD_8.a_inv = "false";
defparam carry_9_5__ADD_8.PCK_LOCATION = "C14R8.lp0.add2.add0";
LUT6 ii2645 (
	. xy ( \ii2645|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2645.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.lut_0";
defparam ii2645.PCK_LOCATION = "C18R11.lp0.lut_0";
defparam ii2645.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[0] .always_en = 1;
LUT6 ii2646 (
	. xy ( \ii2646|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \ii2645|xy_net  ),
	. f2 ( \ii2644|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2643|xy_net  )
);
defparam ii2646.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.lut_0";
defparam ii2646.PCK_LOCATION = "C18R12.lp0.lut_0";
defparam ii2646.config_data = 64'b0101010101010101000011110000001101010101010101010000111100000011;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15]|qx_net  ),
	. di ( \ii2877|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[15] .always_en = 1;
LUT6 ii2647 (
	. xy ( \ii2647|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2647.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2647.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2647.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7]|qx_net  ),
	. di ( \ii2923|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[7] .always_en = 1;
LUT6 ii2648 (
	. xy ( \ii2648|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[10]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2648.PLACE_LOCATION = "C16R8.le_tile.le_guts.lp0.lut_0";
defparam ii2648.PCK_LOCATION = "C16R8.lp0.lut_0";
defparam ii2648.config_data = 64'b0001101100011011000110110001101100011011000110110001101100011011;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[6]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[22] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[3] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[4]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[4] .always_en = 1;
LUT6 ii2649 (
	. xy ( \ii2649|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]|qx_net  ),
	. f2 ( \ii2648|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2649.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2649.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2649.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
LUT6 ii2650 (
	. xy ( \ii2650|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[2]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[18]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[2]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[2]|qx_net  )
);
defparam ii2650.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2650.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2650.config_data = 64'b1100101011111111110010100000111111001010111100001100101000000000;
REG \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9]|qx_net  ),
	. di ( \ii2338|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( \ii2301|xy_net  ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .PLACE_LOCATION = "C10R5.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .PCK_LOCATION = "C10R5.lp0.reg0";
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_sc1_data_cnt_reg[9] .always_en = 0;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. di ( \ii2679|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .PLACE_LOCATION = "C10R11.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .PCK_LOCATION = "C10R11.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23] .always_en = 1;
LUT6 ii2651 (
	. xy ( \ii2651|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2650|xy_net  ),
	. f1 ( \ii2649|xy_net  ),
	. f0 ( \ii2647|xy_net  )
);
defparam ii2651.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2651.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2651.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8]|qx_net  ),
	. di ( \ii3166|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .PLACE_LOCATION = "C20R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .PCK_LOCATION = "C20R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_5_In2p_reg[8] .always_en = 1;
LUT6 ii2652 (
	. xy ( \ii2652|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2652.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2652.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2652.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
LUT6 ii2653 (
	. xy ( \ii2653|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[11]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2653.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2653.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2653.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2654 (
	. xy ( \ii2654|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]|qx_net  ),
	. f2 ( \ii2653|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2654.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2654.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2654.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
REG uut_dataReadBack_mipi_periph_tx_cmd_req_reg (
	. qx ( \uut_dataReadBack_mipi_periph_tx_cmd_req_reg|qx_net  ),
	. di ( \ii3388|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.latch_mode = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.init = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.PLACE_LOCATION = "C4R6.le_tile.le_guts.lp0.reg0";
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.sr_inv = 1;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.sync_mode = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.no_sr = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.sr_value = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.PCK_LOCATION = "C4R6.lp0.reg0";
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.clk_inv = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.en_inv = 0;
defparam uut_dataReadBack_mipi_periph_tx_cmd_req_reg.always_en = 1;
LUT6 ii2655 (
	. xy ( \ii2655|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[3]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[19]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[3]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[3]|qx_net  )
);
defparam ii2655.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2655.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2655.config_data = 64'b1100101011111111110010100000111111001010111100001100101000000000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[1] .always_en = 1;
LUT6 ii2656 (
	. xy ( \ii2656|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2655|xy_net  ),
	. f1 ( \ii2654|xy_net  ),
	. f0 ( \ii2652|xy_net  )
);
defparam ii2656.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2656.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2656.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16]|qx_net  ),
	. di ( \ii2879|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[16] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0]|qx_net  ),
	. di ( \carry_9_13__ADD_0|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[0] .always_en = 1;
LUT6 ii2657 (
	. xy ( \ii2657|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_10_reg[1]|qx_net  )
);
defparam ii2657.PLACE_LOCATION = "C18R12.le_tile.le_guts.lp0.lut_0";
defparam ii2657.PCK_LOCATION = "C18R12.lp0.lut_0";
defparam ii2657.config_data = 64'b1100110010101010111111111111000011001100101010100000000011110000;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[0]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .PCK_LOCATION = "C20R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8]|qx_net  ),
	. di ( \ii2925|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[8] .always_en = 1;
LUT6 ii2658 (
	. xy ( \ii2658|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]|qx_net  ),
	. f1 ( \ii2657|xy_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2658.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2658.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2658.config_data = 64'b0011001100001010000000000000000000110011010111110000000000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[7]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[23] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[8]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .PLACE_LOCATION = "C18R19.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .PCK_LOCATION = "C18R19.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[4] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[5]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[5] .always_en = 1;
LUT6 ii2659 (
	. xy ( \ii2659|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_13_reg[1]|qx_net  ),
	. f2 ( \ii2612|xy_net  ),
	. f1 ( \ii2582|xy_net  ),
	. f0 ( \ii2658|xy_net  )
);
defparam ii2659.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.lut_0";
defparam ii2659.PCK_LOCATION = "C18R11.lp0.lut_0";
defparam ii2659.config_data = 64'b0101010101010101010101010000000101010101010101010101010000000000;
LUT6 ii2660 (
	. xy ( \ii2660|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2660.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2660.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2660.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. di ( \ii2684|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .PLACE_LOCATION = "C10R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .PCK_LOCATION = "C10R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24] .always_en = 1;
LUT6 ii2661 (
	. xy ( \ii2661|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[12]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2661.PLACE_LOCATION = "C16R9.le_tile.le_guts.lp0.lut_0";
defparam ii2661.PCK_LOCATION = "C16R9.lp0.lut_0";
defparam ii2661.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
LUT6 ii2662 (
	. xy ( \ii2662|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]|qx_net  ),
	. f2 ( \ii2661|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2662.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2662.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2662.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
LUT6 ii2663 (
	. xy ( \ii2663|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[4]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[20]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[4]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[4]|qx_net  )
);
defparam ii2663.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2663.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2663.config_data = 64'b1100101011111111110010100000111111001010111100001100101000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[0] .always_en = 1;
LUT6 ii2664 (
	. xy ( \ii2664|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2663|xy_net  ),
	. f1 ( \ii2662|xy_net  ),
	. f0 ( \ii2660|xy_net  )
);
defparam ii2664.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.lut_0";
defparam ii2664.PCK_LOCATION = "C18R11.lp0.lut_0";
defparam ii2664.config_data = 64'b1111000001010101001100110011001111110000010101010011001100110011;
LUT6 ii2665 (
	. xy ( \ii2665|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2665.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2665.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2665.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d1_reg|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.latch_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.init = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.PLACE_LOCATION = "C16R24.le_tile.le_guts.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.sr_inv = 1;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.sync_mode = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.no_sr = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.sr_value = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.PCK_LOCATION = "C16R24.lp0.reg0";
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.clk_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.en_inv = 0;
defparam glue_rx_packet_tx_packet_mipi_tx_packet_generator_mipi_tx_timing_generator_inst_hsync_d2_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[2] .always_en = 1;
LUT6 ii2666 (
	. xy ( \ii2666|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[13]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2666.PLACE_LOCATION = "C18R8.le_tile.le_guts.lp0.lut_0";
defparam ii2666.PCK_LOCATION = "C18R8.lp0.lut_0";
defparam ii2666.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[0]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17]|qx_net  ),
	. di ( \ii2881|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .PLACE_LOCATION = "C6R21.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .PCK_LOCATION = "C6R21.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[17] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1]|qx_net  ),
	. di ( \carry_9_13__ADD_1|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[1] .always_en = 1;
LUT6 ii2667 (
	. xy ( \ii2667|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]|qx_net  ),
	. f2 ( \ii2666|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2667.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2667.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2667.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[1]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .PLACE_LOCATION = "C20R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .PCK_LOCATION = "C20R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9]|qx_net  ),
	. di ( \ii2927|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .PLACE_LOCATION = "C10R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .PCK_LOCATION = "C10R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[9] .always_en = 1;
LUT6 ii2668 (
	. xy ( \ii2668|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[5]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[21]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[5]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[5]|qx_net  )
);
defparam ii2668.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2668.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2668.config_data = 64'b1100101011111111110010100000111111001010111100001100101000000000;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[8]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .PLACE_LOCATION = "C16R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .PCK_LOCATION = "C16R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[24] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5]|qx_net  ),
	. di ( \GND_0_inst|Y_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .PLACE_LOCATION = "C16R17.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .PCK_LOCATION = "C16R17.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_10_In1p_reg[5] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[6]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[6] .always_en = 1;
LUT6 ii2669 (
	. xy ( \ii2669|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2668|xy_net  ),
	. f1 ( \ii2667|xy_net  ),
	. f0 ( \ii2665|xy_net  )
);
defparam ii2669.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2669.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2669.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2670 (
	. xy ( \ii2670|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2670.PLACE_LOCATION = "C18R8.le_tile.le_guts.lp0.lut_0";
defparam ii2670.PCK_LOCATION = "C18R8.lp0.lut_0";
defparam ii2670.config_data = 64'b0010011100100111001001110010011100100111001001110010011100100111;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. di ( \ii2688|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25] .always_en = 1;
LUT6 ii2671 (
	. xy ( \ii2671|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[14]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2671.PLACE_LOCATION = "C16R7.le_tile.le_guts.lp0.lut_0";
defparam ii2671.PCK_LOCATION = "C16R7.lp0.lut_0";
defparam ii2671.config_data = 64'b0001101100011011000110110001101100011011000110110001101100011011;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[19]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[0] .always_en = 1;
LUT6 ii2672 (
	. xy ( \ii2672|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]|qx_net  ),
	. f2 ( \ii2671|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2672.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2672.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2672.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
LUT6 ii2673 (
	. xy ( \ii2673|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[6]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[22]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[6]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[6]|qx_net  )
);
defparam ii2673.PLACE_LOCATION = "C16R11.le_tile.le_guts.lp0.lut_0";
defparam ii2673.PCK_LOCATION = "C16R11.lp0.lut_0";
defparam ii2673.config_data = 64'b1100101011111111110010100000111111001010111100001100101000000000;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[1] .always_en = 1;
LUT6 ii2674 (
	. xy ( \ii2674|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2673|xy_net  ),
	. f1 ( \ii2672|xy_net  ),
	. f0 ( \ii2670|xy_net  )
);
defparam ii2674.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2674.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2674.config_data = 64'b1111000001010101001100110011001111110000010101010011001100110011;
LUT6 ii2675 (
	. xy ( \ii2675|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2675.PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.lut_0";
defparam ii2675.PCK_LOCATION = "C20R8.lp0.lut_0";
defparam ii2675.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .PLACE_LOCATION = "C18R15.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .PCK_LOCATION = "C18R15.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_9_In1p_reg[3] .always_en = 1;
LUT6 ii2676 (
	. xy ( \ii2676|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[15]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2676.PLACE_LOCATION = "C18R8.le_tile.le_guts.lp0.lut_0";
defparam ii2676.PCK_LOCATION = "C18R8.lp0.lut_0";
defparam ii2676.config_data = 64'b0001101100011011000110110001101100011011000110110001101100011011;
REG \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]|qx_net  ),
	. di ( \ii2479|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .PCK_LOCATION = "C16R10.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[1]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .PLACE_LOCATION = "C16R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .PCK_LOCATION = "C16R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t3_out1_1_reg[1] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18]|qx_net  ),
	. di ( \ii2883|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .PLACE_LOCATION = "C8R22.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .PCK_LOCATION = "C8R22.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t83_out1_1_reg[18] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2]|qx_net  ),
	. di ( \carry_9_13__ADD_2|s_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .PLACE_LOCATION = "C16R16.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .PCK_LOCATION = "C16R16.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_11_In2p_reg[2] .always_en = 1;
LUT6 ii2677 (
	. xy ( \ii2677|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]|qx_net  ),
	. f2 ( \ii2676|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2677.PLACE_LOCATION = "C20R9.le_tile.le_guts.lp0.lut_0";
defparam ii2677.PCK_LOCATION = "C20R9.lp0.lut_0";
defparam ii2677.config_data = 64'b1100000011100010110100011111001111000000111000101101000111110011;
REG \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_u_t7_ram_d1|doa[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .PLACE_LOCATION = "C18R14.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .PCK_LOCATION = "C18R14.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t102_out1_reg[2] .always_en = 1;
LUT6 ii2678 (
	. xy ( \ii2678|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[7]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[23]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_7_reg[7]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[7]|qx_net  )
);
defparam ii2678.PLACE_LOCATION = "C18R10.le_tile.le_guts.lp0.lut_0";
defparam ii2678.PCK_LOCATION = "C18R10.lp0.lut_0";
defparam ii2678.config_data = 64'b1100101011111111110010100000111111001010111100001100101000000000;
REG \glue_rx_packet_tx_packet_rx_payload_d_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_rx_payload_d_reg[10]|qx_net  ),
	. di ( \mipi_inst_u_mipi1|periph_rx_payload[10]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .PLACE_LOCATION = "C4R7.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .PCK_LOCATION = "C4R7.lp0.reg0";
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_rx_payload_d_reg[10] .always_en = 1;
REG \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25]  (
	. qx ( \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_from_sc_fifo_u1_hardfifo_u_inst|dout[9]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_gbuf_u_gbuf|out_net  )
);
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .init = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .PLACE_LOCATION = "C14R28.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .PCK_LOCATION = "C14R28.lp0.reg0";
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_mipi_tx_packet_generator_host_tx_payload_reg[25] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t9_out1_9_reg[7]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .PLACE_LOCATION = "C20R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .PCK_LOCATION = "C20R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_6_In3p_reg[7] .always_en = 1;
LUT6 ii2679 (
	. xy ( \ii2679|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2678|xy_net  ),
	. f1 ( \ii2677|xy_net  ),
	. f0 ( \ii2675|xy_net  )
);
defparam ii2679.PLACE_LOCATION = "C18R9.le_tile.le_guts.lp0.lut_0";
defparam ii2679.PCK_LOCATION = "C18R9.lp0.lut_0";
defparam ii2679.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2680 (
	. xy ( \ii2680|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f0 ( \ii2609|xy_net  )
);
defparam ii2680.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2680.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2680.config_data = 64'b1101100011011000110110001101100011011000110110001101100011011000;
REG mcu_arbiter_reg_sel_reg (
	. qx ( \mcu_arbiter_reg_sel_reg|qx_net  ),
	. di ( \ii2038|xy_net  ),
	. sr ( ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO3_net  )
);
defparam mcu_arbiter_reg_sel_reg.latch_mode = 0;
defparam mcu_arbiter_reg_sel_reg.init = 0;
defparam mcu_arbiter_reg_sel_reg.PLACE_LOCATION = "C4R20.le_tile.le_guts.lp0.reg0";
defparam mcu_arbiter_reg_sel_reg.sr_inv = 0;
defparam mcu_arbiter_reg_sel_reg.sync_mode = 1;
defparam mcu_arbiter_reg_sel_reg.no_sr = 1;
defparam mcu_arbiter_reg_sel_reg.sr_value = 0;
defparam mcu_arbiter_reg_sel_reg.PCK_LOCATION = "C4R20.lp0.reg0";
defparam mcu_arbiter_reg_sel_reg.clk_inv = 0;
defparam mcu_arbiter_reg_sel_reg.en_inv = 0;
defparam mcu_arbiter_reg_sel_reg.always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26]|qx_net  ),
	. di ( \ii2693|xy_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .PLACE_LOCATION = "C6R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .PCK_LOCATION = "C6R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[26] .always_en = 1;
LUT6 ii2681 (
	. xy ( \ii2681|xy_net  ),
	. f5 ( ),
	. f4 ( ),
	. f3 ( ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[16]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_reg_2_[1]|qx_net  )
);
defparam ii2681.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2681.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2681.config_data = 64'b1110010011100100111001001110010011100100111001001110010011100100;
REG \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t45_out1_reg[20]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .PLACE_LOCATION = "C8R12.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .sync_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .PCK_LOCATION = "C8R12.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_u_MAC_0_In1p_reg[1] .always_en = 1;
LUT6 ii2682 (
	. xy ( \ii2682|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f2 ( \ii2681|xy_net  ),
	. f1 ( \ii2612|xy_net  ),
	. f0 ( \ii2582|xy_net  )
);
defparam ii2682.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2682.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2682.config_data = 64'b0000110000101110000111010011111100001100001011100001110100111111;
LUT6 ii2683 (
	. xy ( \ii2683|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[8]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[24]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[0]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[0]|qx_net  )
);
defparam ii2683.PLACE_LOCATION = "C18R11.le_tile.le_guts.lp0.lut_0";
defparam ii2683.PCK_LOCATION = "C18R11.lp0.lut_0";
defparam ii2683.config_data = 64'b1011111110001111101100111000001110111100100011001011000010000000;
REG \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_to_sc_fifo_u1_hardfifo_u_inst|dout[2]_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .PLACE_LOCATION = "C10R6.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .PCK_LOCATION = "C10R6.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t10_out1_1_reg[10] .always_en = 1;
REG \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2]  (
	. qx ( \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2]|qx_net  ),
	. di ( \glue_rx_packet_tx_packet_u_scaler_t72_out1_reg[2]|qx_net  ),
	. sr ( \ii1982_dup|xy_net  ),
	. en ( ),
	. clk ( \u_pll_pll_u0|CO0_net  )
);
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .latch_mode = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .init = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .PLACE_LOCATION = "C20R8.le_tile.le_guts.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .sr_inv = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .sync_mode = 1;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .no_sr = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .sr_value = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .PCK_LOCATION = "C20R8.lp0.reg0";
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .clk_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .en_inv = 0;
defparam \glue_rx_packet_tx_packet_u_scaler_t44_out1_1_reg[2] .always_en = 1;
LUT6 ii2684 (
	. xy ( \ii2684|xy_net  ),
	. f5 ( ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[3]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[2]|qx_net  ),
	. f2 ( \ii2683|xy_net  ),
	. f1 ( \ii2682|xy_net  ),
	. f0 ( \ii2680|xy_net  )
);
defparam ii2684.PLACE_LOCATION = "C20R11.le_tile.le_guts.lp0.lut_0";
defparam ii2684.PCK_LOCATION = "C20R11.lp0.lut_0";
defparam ii2684.config_data = 64'b1111000010101010001100110011001111110000101010100011001100110011;
LUT6 ii2685 (
	. xy ( \ii2685|xy_net  ),
	. f5 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[9]|qx_net  ),
	. f4 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[25]|qx_net  ),
	. f3 ( \glue_rx_packet_tx_packet_u_scaler_t52_out1_1_reg[1]|qx_net  ),
	. f2 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[1]|qx_net  ),
	. f1 ( \glue_rx_packet_tx_packet_u_scaler_t35_reg_dul_reg_2_[0]|qx_net  ),
	. f0 ( \glue_rx_packet_tx_packet_u_scaler_t1_out1_4_reg[1]|qx_net  )
);
defparam ii2685.PLACE_LOCATION = "C16R10.le_tile.le_guts.lp0.lut_0";
defparam ii2685.PCK_LOCATION = "C16R10.lp0.lut_0";
defparam ii2685.config_data = 64'b1011111110001111101100111000001110111100100011001011000010000000;
endmodule // mipi_rx_pinf_tx_pinf_1080
